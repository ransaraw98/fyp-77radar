`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 05/23/2023 02:45:31 PM
// Design Name: 
// Module Name: rom
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module sp_rom #(
    parameter integer ADDRW = 14,
    parameter integer DATA_WIDTH = 32,
    parameter RAM_TYPE = "block"
)
(
input [ADDRW-1:0] addr,
input clk,
input en,
output wire [DATA_WIDTH-1:0] dout
    );
    
//DD clock
reg r_clk50=0;

wire w_xor_clk50=(r_clk50 ^ clk);

always@(posedge w_xor_clk50) begin

    r_clk50=~r_clk50;

    // your code on both neg/pos
end
 
    
 (*rom_style = RAM_TYPE*) reg [DATA_WIDTH-1:0] data;   
    
always@(posedge w_xor_clk50)
begin
    if(en)
    case (addr)
        14'd0:data <=32'h0001FFFF;14'd1:data <=32'hFF850027;14'd2:data <=32'hFF370066;
14'd3:data <=32'hFF7500D6;14'd4:data <=32'hFFB700FD;14'd5:data <=32'hFFE900EF;
14'd6:data <=32'h001200D7;14'd7:data <=32'h002C00B0;14'd8:data <=32'h00390091;
14'd9:data <=32'h003D0075;14'd10:data <=32'h003C005D;14'd11:data <=32'h0033004A;
14'd12:data <=32'h0028003C;14'd13:data <=32'h00190035;14'd14:data <=32'h000A0037;
14'd15:data <=32'hFFFE0041;14'd16:data <=32'hFFF80053;14'd17:data <=32'hFFFC0067;
14'd18:data <=32'h000C007A;14'd19:data <=32'h00250086;14'd20:data <=32'h00420088;
14'd21:data <=32'h0061007E;14'd22:data <=32'h0079006A;14'd23:data <=32'h0089004F;
14'd24:data <=32'h00900034;14'd25:data <=32'h008F001B;14'd26:data <=32'h00890004;
14'd27:data <=32'h0080FFF4;14'd28:data <=32'h0076FFE6;14'd29:data <=32'h006AFFDA;
14'd30:data <=32'h005FFFCF;14'd31:data <=32'h0051FFC9;14'd32:data <=32'h0042FFC4;
14'd33:data <=32'h0032FFC4;14'd34:data <=32'h0025FFC9;14'd35:data <=32'h001AFFD0;
14'd36:data <=32'h0013FFDA;14'd37:data <=32'h0012FFE4;14'd38:data <=32'h0014FFED;
14'd39:data <=32'h0018FFF4;14'd40:data <=32'h001EFFF7;14'd41:data <=32'h0021FFFA;
14'd42:data <=32'h0026FFFE;14'd43:data <=32'h002A0003;14'd44:data <=32'h00340008;
14'd45:data <=32'h0043000D;14'd46:data <=32'h0058000C;14'd47:data <=32'h00720003;
14'd48:data <=32'h008CFFF0;14'd49:data <=32'h00A1FFCF;14'd50:data <=32'h00ACFFA6;
14'd51:data <=32'h00ABFF77;14'd52:data <=32'h009CFF46;14'd53:data <=32'h007EFF19;
14'd54:data <=32'h0055FEF3;14'd55:data <=32'h0021FED9;14'd56:data <=32'hFFE8FEC9;
14'd57:data <=32'hFFABFEC6;14'd58:data <=32'hFF6CFED1;14'd59:data <=32'hFF2EFEEB;
14'd60:data <=32'hFEF6FF12;14'd61:data <=32'hFEC7FF4A;14'd62:data <=32'hFEA6FF8D;
14'd63:data <=32'hFE98FFD8;14'd64:data <=32'hFF5EFFAB;14'd65:data <=32'hFF39FFBD;
14'd66:data <=32'hFF0DFFCF;14'd67:data <=32'hFEBE0007;14'd68:data <=32'hFF080065;
14'd69:data <=32'hFF2B007D;14'd70:data <=32'hFF4B008C;14'd71:data <=32'hFF6A0094;
14'd72:data <=32'hFF830098;14'd73:data <=32'hFF9A009D;14'd74:data <=32'hFFB0009D;
14'd75:data <=32'hFFC6009C;14'd76:data <=32'hFFD80096;14'd77:data <=32'hFFE8008E;
14'd78:data <=32'hFFF30086;14'd79:data <=32'hFFFB0080;14'd80:data <=32'h0001007C;
14'd81:data <=32'h0009007B;14'd82:data <=32'h0014007B;14'd83:data <=32'h00230078;
14'd84:data <=32'h00340072;14'd85:data <=32'h00420064;14'd86:data <=32'h004B0053;
14'd87:data <=32'h004D003D;14'd88:data <=32'h0048002B;14'd89:data <=32'h003C0020;
14'd90:data <=32'h002F001A;14'd91:data <=32'h0024001E;14'd92:data <=32'h001E0025;
14'd93:data <=32'h001E002E;14'd94:data <=32'h00240035;14'd95:data <=32'h002B0039;
14'd96:data <=32'h00350039;14'd97:data <=32'h00400035;14'd98:data <=32'h00470030;
14'd99:data <=32'h004D0028;14'd100:data <=32'h0053001F;14'd101:data <=32'h00570015;
14'd102:data <=32'h00590009;14'd103:data <=32'h0056FFFD;14'd104:data <=32'h0050FFF2;
14'd105:data <=32'h0046FFE9;14'd106:data <=32'h0038FFE6;14'd107:data <=32'h002AFFEA;
14'd108:data <=32'h001FFFF5;14'd109:data <=32'h001B0006;14'd110:data <=32'h0021001B;
14'd111:data <=32'h0032002C;14'd112:data <=32'h004D0037;14'd113:data <=32'h006E0035;
14'd114:data <=32'h00900027;14'd115:data <=32'h00AE000C;14'd116:data <=32'h00C3FFE7;
14'd117:data <=32'h00CCFFBD;14'd118:data <=32'h00C9FF8E;14'd119:data <=32'h00BCFF63;
14'd120:data <=32'h00A5FF39;14'd121:data <=32'h0086FF14;14'd122:data <=32'h005EFEF7;
14'd123:data <=32'h002FFEE0;14'd124:data <=32'hFFF9FED5;14'd125:data <=32'hFFC0FED7;
14'd126:data <=32'hFF88FEE7;14'd127:data <=32'hFF57FF05;14'd128:data <=32'hFF73FEF8;
14'd129:data <=32'hFF36FF09;14'd130:data <=32'hFF14FF1E;14'd131:data <=32'hFF57FF1F;
14'd132:data <=32'hFF71FF66;14'd133:data <=32'hFF63FF71;14'd134:data <=32'hFF51FF7D;
14'd135:data <=32'hFF3CFF8C;14'd136:data <=32'hFF26FFA3;14'd137:data <=32'hFF11FFC2;
14'd138:data <=32'hFF04FFE9;14'd139:data <=32'hFF020013;14'd140:data <=32'hFF08003E;
14'd141:data <=32'hFF180065;14'd142:data <=32'hFF2E0088;14'd143:data <=32'hFF4B00A7;
14'd144:data <=32'hFF6C00BF;14'd145:data <=32'hFF9300D0;14'd146:data <=32'hFFBD00DB;
14'd147:data <=32'hFFEA00DB;14'd148:data <=32'h001700CF;14'd149:data <=32'h003F00B6;
14'd150:data <=32'h005C0093;14'd151:data <=32'h006D006A;14'd152:data <=32'h006E003E;
14'd153:data <=32'h00620018;14'd154:data <=32'h0049FFFD;14'd155:data <=32'h002DFFEF;
14'd156:data <=32'h000FFFEC;14'd157:data <=32'hFFF8FFF3;14'd158:data <=32'hFFE50002;
14'd159:data <=32'hFFDB0013;14'd160:data <=32'hFFD70025;14'd161:data <=32'hFFD80037;
14'd162:data <=32'hFFDE0048;14'd163:data <=32'hFFE80056;14'd164:data <=32'hFFF50062;
14'd165:data <=32'h0006006B;14'd166:data <=32'h0019006E;14'd167:data <=32'h002C006C;
14'd168:data <=32'h003C0064;14'd169:data <=32'h004A0057;14'd170:data <=32'h0052004B;
14'd171:data <=32'h0055003F;14'd172:data <=32'h00520037;14'd173:data <=32'h00510036;
14'd174:data <=32'h00530037;14'd175:data <=32'h005A003A;14'd176:data <=32'h0067003C;
14'd177:data <=32'h00780038;14'd178:data <=32'h008B002D;14'd179:data <=32'h009C001A;
14'd180:data <=32'h00A60003;14'd181:data <=32'h00ABFFE7;14'd182:data <=32'h00A8FFCF;
14'd183:data <=32'h00A0FFB6;14'd184:data <=32'h0095FFA3;14'd185:data <=32'h0088FF93;
14'd186:data <=32'h007AFF83;14'd187:data <=32'h006CFF76;14'd188:data <=32'h005BFF6A;
14'd189:data <=32'h004AFF60;14'd190:data <=32'h0036FF5A;14'd191:data <=32'h0023FF59;
14'd192:data <=32'h0069FECF;14'd193:data <=32'h002BFEAD;14'd194:data <=32'hFFF2FEB6;
14'd195:data <=32'h0021FF55;14'd196:data <=32'h004BFF7A;14'd197:data <=32'h0046FF5C;
14'd198:data <=32'h0036FF3B;14'd199:data <=32'h001AFF1C;14'd200:data <=32'hFFECFF05;
14'd201:data <=32'hFFB8FEFE;14'd202:data <=32'hFF81FF05;14'd203:data <=32'hFF4EFF1C;
14'd204:data <=32'hFF21FF41;14'd205:data <=32'hFEFFFF6E;14'd206:data <=32'hFEE9FFA0;
14'd207:data <=32'hFEDEFFD5;14'd208:data <=32'hFEDE000E;14'd209:data <=32'hFEEB0045;
14'd210:data <=32'hFF060078;14'd211:data <=32'hFF2C00A3;14'd212:data <=32'hFF5D00C3;
14'd213:data <=32'hFF9400D2;14'd214:data <=32'hFFCC00D1;14'd215:data <=32'hFFFD00BE;
14'd216:data <=32'h002200A1;14'd217:data <=32'h003A007E;14'd218:data <=32'h00430059;
14'd219:data <=32'h00410039;14'd220:data <=32'h0039001F;14'd221:data <=32'h002B000B;
14'd222:data <=32'h001DFFFF;14'd223:data <=32'h000DFFF6;14'd224:data <=32'hFFFDFFF1;
14'd225:data <=32'hFFEEFFEF;14'd226:data <=32'hFFDBFFF1;14'd227:data <=32'hFFCAFFF8;
14'd228:data <=32'hFFBA0004;14'd229:data <=32'hFFAF0016;14'd230:data <=32'hFFA7002B;
14'd231:data <=32'hFFA60041;14'd232:data <=32'hFFAA0058;14'd233:data <=32'hFFB4006D;
14'd234:data <=32'hFFC00080;14'd235:data <=32'hFFCF0091;14'd236:data <=32'hFFE200A1;
14'd237:data <=32'hFFF700B0;14'd238:data <=32'h001300BC;14'd239:data <=32'h003300C4;
14'd240:data <=32'h005A00C6;14'd241:data <=32'h008400BD;14'd242:data <=32'h00AC00A7;
14'd243:data <=32'h00CD0085;14'd244:data <=32'h00E5005A;14'd245:data <=32'h00EE002A;
14'd246:data <=32'h00EBFFFB;14'd247:data <=32'h00DBFFD3;14'd248:data <=32'h00C2FFB2;
14'd249:data <=32'h00A7FF9D;14'd250:data <=32'h008AFF90;14'd251:data <=32'h006FFF8C;
14'd252:data <=32'h0057FF8D;14'd253:data <=32'h0044FF94;14'd254:data <=32'h0035FF9D;
14'd255:data <=32'h002AFFAA;14'd256:data <=32'h00CCFF9D;14'd257:data <=32'h00C7FF70;
14'd258:data <=32'h009FFF4F;14'd259:data <=32'h0030FF99;14'd260:data <=32'h0066FFCF;
14'd261:data <=32'h0078FFBC;14'd262:data <=32'h0082FF9E;14'd263:data <=32'h0082FF7B;
14'd264:data <=32'h0072FF56;14'd265:data <=32'h0056FF37;14'd266:data <=32'h0031FF22;
14'd267:data <=32'h0006FF17;14'd268:data <=32'hFFDDFF17;14'd269:data <=32'hFFB5FF21;
14'd270:data <=32'hFF93FF31;14'd271:data <=32'hFF73FF47;14'd272:data <=32'hFF59FF64;
14'd273:data <=32'hFF43FF84;14'd274:data <=32'hFF34FFA9;14'd275:data <=32'hFF30FFD1;
14'd276:data <=32'hFF36FFF9;14'd277:data <=32'hFF45001B;14'd278:data <=32'hFF5C0036;
14'd279:data <=32'hFF770046;14'd280:data <=32'hFF90004F;14'd281:data <=32'hFFA60050;
14'd282:data <=32'hFFB7004F;14'd283:data <=32'hFFC5004D;14'd284:data <=32'hFFCF004C;
14'd285:data <=32'hFFDB004B;14'd286:data <=32'hFFE90048;14'd287:data <=32'hFFF70043;
14'd288:data <=32'h00060038;14'd289:data <=32'h00120027;14'd290:data <=32'h00160012;
14'd291:data <=32'h0013FFFB;14'd292:data <=32'h0006FFE7;14'd293:data <=32'hFFF3FFD8;
14'd294:data <=32'hFFDBFFD0;14'd295:data <=32'hFFC1FFCF;14'd296:data <=32'hFFA6FFD6;
14'd297:data <=32'hFF8CFFE5;14'd298:data <=32'hFF76FFFA;14'd299:data <=32'hFF630017;
14'd300:data <=32'hFF58003A;14'd301:data <=32'hFF530063;14'd302:data <=32'hFF590090;
14'd303:data <=32'hFF6E00BE;14'd304:data <=32'hFF9100E7;14'd305:data <=32'hFFC00108;
14'd306:data <=32'hFFF9011A;14'd307:data <=32'h0036011A;14'd308:data <=32'h006F0108;
14'd309:data <=32'h00A000E9;14'd310:data <=32'h00C500BF;14'd311:data <=32'h00DB0092;
14'd312:data <=32'h00E30064;14'd313:data <=32'h00E3003B;14'd314:data <=32'h00DA0017;
14'd315:data <=32'h00CDFFFA;14'd316:data <=32'h00BDFFE2;14'd317:data <=32'h00ABFFCF;
14'd318:data <=32'h0097FFC3;14'd319:data <=32'h0084FFBC;14'd320:data <=32'h006EFFEF;
14'd321:data <=32'h0075FFEC;14'd322:data <=32'h007FFFD8;14'd323:data <=32'h0092FF97;
14'd324:data <=32'h00B1FFC4;14'd325:data <=32'h00B1FFAE;14'd326:data <=32'h00ABFF95;
14'd327:data <=32'h00A0FF79;14'd328:data <=32'h008AFF5D;14'd329:data <=32'h006BFF49;
14'd330:data <=32'h0046FF3D;14'd331:data <=32'h0022FF3E;14'd332:data <=32'h0002FF47;
14'd333:data <=32'hFFE9FF57;14'd334:data <=32'hFFD8FF69;14'd335:data <=32'hFFCDFF7B;
14'd336:data <=32'hFFC6FF8A;14'd337:data <=32'hFFC2FF98;14'd338:data <=32'hFFBFFFA4;
14'd339:data <=32'hFFBEFFAF;14'd340:data <=32'hFFBEFFBA;14'd341:data <=32'hFFC2FFC0;
14'd342:data <=32'hFFC6FFC5;14'd343:data <=32'hFFCAFFC5;14'd344:data <=32'hFFC9FFC1;
14'd345:data <=32'hFFC1FFBD;14'd346:data <=32'hFFB7FFBB;14'd347:data <=32'hFFA7FFBF;
14'd348:data <=32'hFF97FFCD;14'd349:data <=32'hFF8CFFE1;14'd350:data <=32'hFF89FFF7;
14'd351:data <=32'hFF910010;14'd352:data <=32'hFFA00024;14'd353:data <=32'hFFB60031;
14'd354:data <=32'hFFCD0035;14'd355:data <=32'hFFE3002E;14'd356:data <=32'hFFF30021;
14'd357:data <=32'hFFFD000F;14'd358:data <=32'hFFFEFFFB;14'd359:data <=32'hFFFAFFE8;
14'd360:data <=32'hFFEFFFD7;14'd361:data <=32'hFFDFFFCB;14'd362:data <=32'hFFC8FFC1;
14'd363:data <=32'hFFAFFFBE;14'd364:data <=32'hFF92FFC4;14'd365:data <=32'hFF75FFD2;
14'd366:data <=32'hFF5BFFEB;14'd367:data <=32'hFF46000D;14'd368:data <=32'hFF3D0036;
14'd369:data <=32'hFF410062;14'd370:data <=32'hFF51008B;14'd371:data <=32'hFF6C00AD;
14'd372:data <=32'hFF8D00C6;14'd373:data <=32'hFFB000D5;14'd374:data <=32'hFFD100DC;
14'd375:data <=32'hFFEF00DB;14'd376:data <=32'h000900DA;14'd377:data <=32'h002200D8;
14'd378:data <=32'h003A00D5;14'd379:data <=32'h005400D0;14'd380:data <=32'h007000C9;
14'd381:data <=32'h008C00BC;14'd382:data <=32'h00A700AB;14'd383:data <=32'h00BE0094;
14'd384:data <=32'h0080FFF7;14'd385:data <=32'h0075FFF8;14'd386:data <=32'h0078000B;
14'd387:data <=32'h00ED0065;14'd388:data <=32'h01280077;14'd389:data <=32'h013D003F;
14'd390:data <=32'h01450001;14'd391:data <=32'h0140FFC3;14'd392:data <=32'h0128FF83;
14'd393:data <=32'h00FFFF4E;14'd394:data <=32'h00C9FF27;14'd395:data <=32'h008CFF14;
14'd396:data <=32'h0051FF12;14'd397:data <=32'h001DFF20;14'd398:data <=32'hFFF5FF3A;
14'd399:data <=32'hFFD9FF5A;14'd400:data <=32'hFFC8FF7A;14'd401:data <=32'hFFC1FF98;
14'd402:data <=32'hFFC2FFB4;14'd403:data <=32'hFFC8FFCC;14'd404:data <=32'hFFD5FFDF;
14'd405:data <=32'hFFE7FFED;14'd406:data <=32'hFFFAFFF0;14'd407:data <=32'h000DFFEC;
14'd408:data <=32'h001EFFDF;14'd409:data <=32'h0025FFCC;14'd410:data <=32'h0023FFB6;
14'd411:data <=32'h0017FFA3;14'd412:data <=32'h0004FF97;14'd413:data <=32'hFFEEFF92;
14'd414:data <=32'hFFD8FF98;14'd415:data <=32'hFFC6FFA4;14'd416:data <=32'hFFBEFFB4;
14'd417:data <=32'hFFBAFFC3;14'd418:data <=32'hFFBBFFCF;14'd419:data <=32'hFFC0FFD7;
14'd420:data <=32'hFFC3FFDA;14'd421:data <=32'hFFC7FFDD;14'd422:data <=32'hFFC7FFDC;
14'd423:data <=32'hFFC6FFDD;14'd424:data <=32'hFFC5FFDE;14'd425:data <=32'hFFC4FFDF;
14'd426:data <=32'hFFC3FFDE;14'd427:data <=32'hFFBFFFDE;14'd428:data <=32'hFFBCFFDC;
14'd429:data <=32'hFFB4FFDB;14'd430:data <=32'hFFAAFFDD;14'd431:data <=32'hFFA0FFE2;
14'd432:data <=32'hFF96FFEB;14'd433:data <=32'hFF8FFFF6;14'd434:data <=32'hFF8C0002;
14'd435:data <=32'hFF8B000B;14'd436:data <=32'hFF8B0014;14'd437:data <=32'hFF890018;
14'd438:data <=32'hFF81001E;14'd439:data <=32'hFF760027;14'd440:data <=32'hFF670035;
14'd441:data <=32'hFF59004F;14'd442:data <=32'hFF500071;14'd443:data <=32'hFF51009A;
14'd444:data <=32'hFF6000C7;14'd445:data <=32'hFF7C00F2;14'd446:data <=32'hFFA50116;
14'd447:data <=32'hFFD6012F;14'd448:data <=32'h0055008B;14'd449:data <=32'h0059008B;
14'd450:data <=32'h004C0098;14'd451:data <=32'h001E011E;14'd452:data <=32'h007E0154;
14'd453:data <=32'h00C20138;14'd454:data <=32'h00FE010B;14'd455:data <=32'h012D00D0;
14'd456:data <=32'h014B0088;14'd457:data <=32'h0153003D;14'd458:data <=32'h0146FFF6;
14'd459:data <=32'h0127FFB9;14'd460:data <=32'h00FEFF8C;14'd461:data <=32'h00CFFF6F;
14'd462:data <=32'h00A1FF5F;14'd463:data <=32'h0078FF5B;14'd464:data <=32'h0054FF5E;
14'd465:data <=32'h0036FF68;14'd466:data <=32'h001BFF74;14'd467:data <=32'h0006FF84;
14'd468:data <=32'hFFF6FF97;14'd469:data <=32'hFFEDFFAC;14'd470:data <=32'hFFEDFFC2;
14'd471:data <=32'hFFF1FFD3;14'd472:data <=32'hFFFBFFDF;14'd473:data <=32'h0007FFE3;
14'd474:data <=32'h0011FFE2;14'd475:data <=32'h0017FFDD;14'd476:data <=32'h0018FFD9;
14'd477:data <=32'h0018FFD5;14'd478:data <=32'h0016FFD4;14'd479:data <=32'h0017FFD5;
14'd480:data <=32'h001CFFD5;14'd481:data <=32'h0022FFD1;14'd482:data <=32'h0029FFCA;
14'd483:data <=32'h002DFFBC;14'd484:data <=32'h002BFFAB;14'd485:data <=32'h0023FF98;
14'd486:data <=32'h0013FF89;14'd487:data <=32'hFFFFFF7E;14'd488:data <=32'hFFE7FF7A;
14'd489:data <=32'hFFD0FF7E;14'd490:data <=32'hFFBAFF87;14'd491:data <=32'hFFA9FF95;
14'd492:data <=32'hFF9DFFA4;14'd493:data <=32'hFF94FFB5;14'd494:data <=32'hFF8EFFC8;
14'd495:data <=32'hFF8DFFD9;14'd496:data <=32'hFF91FFEA;14'd497:data <=32'hFF9AFFF8;
14'd498:data <=32'hFFA60002;14'd499:data <=32'hFFB50004;14'd500:data <=32'hFFC2FFFF;
14'd501:data <=32'hFFCBFFF2;14'd502:data <=32'hFFCAFFDF;14'd503:data <=32'hFFBEFFCB;
14'd504:data <=32'hFFA5FFBD;14'd505:data <=32'hFF83FFBA;14'd506:data <=32'hFF5EFFC4;
14'd507:data <=32'hFF39FFDD;14'd508:data <=32'hFF1D0005;14'd509:data <=32'hFF0D0035;
14'd510:data <=32'hFF0B0069;14'd511:data <=32'hFF16009E;14'd512:data <=32'hFF6B007F;
14'd513:data <=32'hFF6800A8;14'd514:data <=32'hFF6900BC;14'd515:data <=32'hFF5500A9;
14'd516:data <=32'hFF960106;14'd517:data <=32'hFFC60118;14'd518:data <=32'hFFF9011D;
14'd519:data <=32'h002E0116;14'd520:data <=32'h005D0101;14'd521:data <=32'h008300E2;
14'd522:data <=32'h009C00BE;14'd523:data <=32'h00AA009B;14'd524:data <=32'h00B0007A;
14'd525:data <=32'h00B20060;14'd526:data <=32'h00B1004B;14'd527:data <=32'h00B20038;
14'd528:data <=32'h00B30024;14'd529:data <=32'h00B5000D;14'd530:data <=32'h00B2FFF4;
14'd531:data <=32'h00AAFFDB;14'd532:data <=32'h009CFFC4;14'd533:data <=32'h0089FFB2;
14'd534:data <=32'h0073FFA4;14'd535:data <=32'h005DFF9D;14'd536:data <=32'h0048FF99;
14'd537:data <=32'h0034FF99;14'd538:data <=32'h0020FF9C;14'd539:data <=32'h000DFFA3;
14'd540:data <=32'hFFFBFFAE;14'd541:data <=32'hFFEBFFC0;14'd542:data <=32'hFFE3FFD7;
14'd543:data <=32'hFFE3FFF0;14'd544:data <=32'hFFEE0009;14'd545:data <=32'h0002001D;
14'd546:data <=32'h001E0027;14'd547:data <=32'h003D0025;14'd548:data <=32'h00590016;
14'd549:data <=32'h006FFFFE;14'd550:data <=32'h007BFFDE;14'd551:data <=32'h007CFFBD;
14'd552:data <=32'h0073FF9F;14'd553:data <=32'h0062FF85;14'd554:data <=32'h004BFF6F;
14'd555:data <=32'h0032FF62;14'd556:data <=32'h0016FF5B;14'd557:data <=32'hFFFCFF59;
14'd558:data <=32'hFFE2FF5C;14'd559:data <=32'hFFC9FF66;14'd560:data <=32'hFFB5FF75;
14'd561:data <=32'hFFA6FF87;14'd562:data <=32'hFF9DFF9A;14'd563:data <=32'hFF9CFFAC;
14'd564:data <=32'hFFA0FFB9;14'd565:data <=32'hFFA7FFBF;14'd566:data <=32'hFFACFFBE;
14'd567:data <=32'hFFAAFFB7;14'd568:data <=32'hFFA1FFB0;14'd569:data <=32'hFF8FFFA9;
14'd570:data <=32'hFF78FFAC;14'd571:data <=32'hFF5EFFB8;14'd572:data <=32'hFF47FFCE;
14'd573:data <=32'hFF37FFEC;14'd574:data <=32'hFF2F000D;14'd575:data <=32'hFF30002D;
14'd576:data <=32'hFF3EFF99;14'd577:data <=32'hFF04FFBE;14'd578:data <=32'hFEEDFFF1;
14'd579:data <=32'hFF61003E;14'd580:data <=32'hFF8B008B;14'd581:data <=32'hFFA20092;
14'd582:data <=32'hFFB80092;14'd583:data <=32'hFFCC0090;14'd584:data <=32'hFFDC0089;
14'd585:data <=32'hFFE8007E;14'd586:data <=32'hFFEB0076;14'd587:data <=32'hFFE9006F;
14'd588:data <=32'hFFE40073;14'd589:data <=32'hFFE2007E;14'd590:data <=32'hFFE50090;
14'd591:data <=32'hFFF500A4;14'd592:data <=32'h000E00B4;14'd593:data <=32'h002F00BC;
14'd594:data <=32'h005400B8;14'd595:data <=32'h007700A9;14'd596:data <=32'h00950091;
14'd597:data <=32'h00AC0071;14'd598:data <=32'h00BA004E;14'd599:data <=32'h00BF002B;
14'd600:data <=32'h00BD0007;14'd601:data <=32'h00B3FFE3;14'd602:data <=32'h00A0FFC5;
14'd603:data <=32'h0087FFAA;14'd604:data <=32'h0066FF98;14'd605:data <=32'h0041FF92;
14'd606:data <=32'h001CFF97;14'd607:data <=32'hFFFDFFA8;14'd608:data <=32'hFFE6FFC3;
14'd609:data <=32'hFFDCFFE5;14'd610:data <=32'hFFE00004;14'd611:data <=32'hFFEE001F;
14'd612:data <=32'h00040030;14'd613:data <=32'h001D0039;14'd614:data <=32'h00380038;
14'd615:data <=32'h004D0031;14'd616:data <=32'h00600024;14'd617:data <=32'h006E0015;
14'd618:data <=32'h00780005;14'd619:data <=32'h0082FFF2;14'd620:data <=32'h0089FFDF;
14'd621:data <=32'h008DFFC8;14'd622:data <=32'h008CFFAF;14'd623:data <=32'h0086FF95;
14'd624:data <=32'h007BFF7C;14'd625:data <=32'h006AFF66;14'd626:data <=32'h0056FF53;
14'd627:data <=32'h0040FF45;14'd628:data <=32'h0028FF38;14'd629:data <=32'h0011FF2E;
14'd630:data <=32'hFFF6FF23;14'd631:data <=32'hFFD6FF1B;14'd632:data <=32'hFFB1FF19;
14'd633:data <=32'hFF87FF1D;14'd634:data <=32'hFF5BFF2D;14'd635:data <=32'hFF32FF4B;
14'd636:data <=32'hFF10FF74;14'd637:data <=32'hFEFCFFA5;14'd638:data <=32'hFEF5FFDA;
14'd639:data <=32'hFEFD000B;14'd640:data <=32'hFFC8FF58;14'd641:data <=32'hFF8BFF4B;
14'd642:data <=32'hFF47FF62;14'd643:data <=32'hFF250026;14'd644:data <=32'hFF5B007C;
14'd645:data <=32'hFF810086;14'd646:data <=32'hFFA20085;14'd647:data <=32'hFFC0007C;
14'd648:data <=32'hFFD8006A;14'd649:data <=32'hFFE70054;14'd650:data <=32'hFFEA003C;
14'd651:data <=32'hFFE00029;14'd652:data <=32'hFFCD001C;14'd653:data <=32'hFFB6001E;
14'd654:data <=32'hFFA1002D;14'd655:data <=32'hFF960046;14'd656:data <=32'hFF950064;
14'd657:data <=32'hFFA00082;14'd658:data <=32'hFFB7009C;14'd659:data <=32'hFFD400AC;
14'd660:data <=32'hFFF300B3;14'd661:data <=32'h001100B3;14'd662:data <=32'h002F00AB;
14'd663:data <=32'h0049009E;14'd664:data <=32'h0061008D;14'd665:data <=32'h00750077;
14'd666:data <=32'h0083005E;14'd667:data <=32'h008A0041;14'd668:data <=32'h00890023;
14'd669:data <=32'h007F0007;14'd670:data <=32'h006FFFF1;14'd671:data <=32'h005AFFE3;
14'd672:data <=32'h0042FFDE;14'd673:data <=32'h0030FFE1;14'd674:data <=32'h0022FFE8;
14'd675:data <=32'h0019FFF2;14'd676:data <=32'h0015FFFC;14'd677:data <=32'h00130002;
14'd678:data <=32'h00110008;14'd679:data <=32'h0010000E;14'd680:data <=32'h000E0015;
14'd681:data <=32'h000D0022;14'd682:data <=32'h00110030;14'd683:data <=32'h001A0041;
14'd684:data <=32'h002C004F;14'd685:data <=32'h00460059;14'd686:data <=32'h0064005C;
14'd687:data <=32'h00860054;14'd688:data <=32'h00A70043;14'd689:data <=32'h00C40027;
14'd690:data <=32'h00D90005;14'd691:data <=32'h00E9FFDC;14'd692:data <=32'h00F2FFAF;
14'd693:data <=32'h00F0FF7C;14'd694:data <=32'h00E3FF48;14'd695:data <=32'h00C8FF13;
14'd696:data <=32'h009FFEE1;14'd697:data <=32'h0066FEBA;14'd698:data <=32'h0022FEA1;
14'd699:data <=32'hFFD8FE9C;14'd700:data <=32'hFF8DFEAC;14'd701:data <=32'hFF4BFED1;
14'd702:data <=32'hFF18FF05;14'd703:data <=32'hFEF7FF41;14'd704:data <=32'hFFD1FF68;
14'd705:data <=32'hFFB1FF54;14'd706:data <=32'hFF7DFF41;14'd707:data <=32'hFF04FF59;
14'd708:data <=32'hFF17FFC6;14'd709:data <=32'hFF23FFEB;14'd710:data <=32'hFF330009;
14'd711:data <=32'hFF470021;14'd712:data <=32'hFF5E0032;14'd713:data <=32'hFF760039;
14'd714:data <=32'hFF88003A;14'd715:data <=32'hFF940036;14'd716:data <=32'hFF980031;
14'd717:data <=32'hFF970031;14'd718:data <=32'hFF930037;14'd719:data <=32'hFF920043;
14'd720:data <=32'hFF960054;14'd721:data <=32'hFFA20063;14'd722:data <=32'hFFB30070;
14'd723:data <=32'hFFC60074;14'd724:data <=32'hFFD90074;14'd725:data <=32'hFFE9006F;
14'd726:data <=32'hFFF40066;14'd727:data <=32'hFFFB005F;14'd728:data <=32'hFFFF005A;
14'd729:data <=32'h00040055;14'd730:data <=32'h00080053;14'd731:data <=32'h000C0050;
14'd732:data <=32'h000F004C;14'd733:data <=32'h00130048;14'd734:data <=32'h00140045;
14'd735:data <=32'h00150045;14'd736:data <=32'h00160045;14'd737:data <=32'h001A0047;
14'd738:data <=32'h00220049;14'd739:data <=32'h002C0048;14'd740:data <=32'h00380040;
14'd741:data <=32'h00410035;14'd742:data <=32'h00440026;14'd743:data <=32'h003F0016;
14'd744:data <=32'h00330009;14'd745:data <=32'h00230001;14'd746:data <=32'h000F0005;
14'd747:data <=32'hFFFF0011;14'd748:data <=32'hFFF50026;14'd749:data <=32'hFFF30040;
14'd750:data <=32'hFFFD0059;14'd751:data <=32'h00110071;14'd752:data <=32'h002D0081;
14'd753:data <=32'h004E008A;14'd754:data <=32'h0074008B;14'd755:data <=32'h009A0081;
14'd756:data <=32'h00C2006D;14'd757:data <=32'h00E5004F;14'd758:data <=32'h01040027;
14'd759:data <=32'h0119FFF3;14'd760:data <=32'h0121FFB8;14'd761:data <=32'h0118FF7A;
14'd762:data <=32'h00FDFF3F;14'd763:data <=32'h00D3FF0D;14'd764:data <=32'h009EFEE9;
14'd765:data <=32'h0063FED6;14'd766:data <=32'h002AFED2;14'd767:data <=32'hFFF6FEDD;
14'd768:data <=32'h0013FEFB;14'd769:data <=32'hFFE8FEE9;14'd770:data <=32'hFFCDFEDC;
14'd771:data <=32'hFFF9FED6;14'd772:data <=32'hFFEAFF18;14'd773:data <=32'hFFCCFF1B;
14'd774:data <=32'hFFAFFF21;14'd775:data <=32'hFF8EFF2D;14'd776:data <=32'hFF73FF3F;
14'd777:data <=32'hFF5BFF55;14'd778:data <=32'hFF46FF6C;14'd779:data <=32'hFF33FF86;
14'd780:data <=32'hFF22FFA4;14'd781:data <=32'hFF15FFC7;14'd782:data <=32'hFF0EFFEE;
14'd783:data <=32'hFF0F001A;14'd784:data <=32'hFF1E0047;14'd785:data <=32'hFF380071;
14'd786:data <=32'hFF5E008F;14'd787:data <=32'hFF8B00A1;14'd788:data <=32'hFFB900A2;
14'd789:data <=32'hFFE10097;14'd790:data <=32'h00000081;14'd791:data <=32'h00130066;
14'd792:data <=32'h001D004B;14'd793:data <=32'h001D0033;14'd794:data <=32'h0017001E;
14'd795:data <=32'h000D000E;14'd796:data <=32'hFFFF0002;14'd797:data <=32'hFFEEFFFC;
14'd798:data <=32'hFFDDFFFD;14'd799:data <=32'hFFCA0003;14'd800:data <=32'hFFBC0010;
14'd801:data <=32'hFFB40023;14'd802:data <=32'hFFB30039;14'd803:data <=32'hFFBB004F;
14'd804:data <=32'hFFC9005F;14'd805:data <=32'hFFDD006A;14'd806:data <=32'hFFF1006B;
14'd807:data <=32'h00030066;14'd808:data <=32'h000D005C;14'd809:data <=32'h00120051;
14'd810:data <=32'h00110049;14'd811:data <=32'h000B0048;14'd812:data <=32'h0007004B;
14'd813:data <=32'h00050053;14'd814:data <=32'h0008005E;14'd815:data <=32'h0012006A;
14'd816:data <=32'h001F0071;14'd817:data <=32'h002F0077;14'd818:data <=32'h00410079;
14'd819:data <=32'h00530078;14'd820:data <=32'h00670074;14'd821:data <=32'h007B006D;
14'd822:data <=32'h00910061;14'd823:data <=32'h00A60051;14'd824:data <=32'h00B70039;
14'd825:data <=32'h00C3001C;14'd826:data <=32'h00C8FFFE;14'd827:data <=32'h00C3FFDF;
14'd828:data <=32'h00B8FFC5;14'd829:data <=32'h00AAFFB3;14'd830:data <=32'h009DFFA6;
14'd831:data <=32'h0094FF9C;14'd832:data <=32'h00ECFF3B;14'd833:data <=32'h00D0FF06;
14'd834:data <=32'h00ABFEF3;14'd835:data <=32'h00B1FF82;14'd836:data <=32'h00C4FFA4;
14'd837:data <=32'h00C3FF7A;14'd838:data <=32'h00B6FF50;14'd839:data <=32'h009CFF26;
14'd840:data <=32'h0079FF04;14'd841:data <=32'h004EFEEA;14'd842:data <=32'h001CFED9;
14'd843:data <=32'hFFE7FED0;14'd844:data <=32'hFFADFED4;14'd845:data <=32'hFF72FEE6;
14'd846:data <=32'hFF3CFF07;14'd847:data <=32'hFF0EFF38;14'd848:data <=32'hFEF0FF74;
14'd849:data <=32'hFEE3FFB6;14'd850:data <=32'hFEECFFF8;14'd851:data <=32'hFF050031;
14'd852:data <=32'hFF2B005C;14'd853:data <=32'hFF580077;14'd854:data <=32'hFF850084;
14'd855:data <=32'hFFAF0084;14'd856:data <=32'hFFD2007A;14'd857:data <=32'hFFEF006B;
14'd858:data <=32'h00040056;14'd859:data <=32'h00120040;14'd860:data <=32'h001B0028;
14'd861:data <=32'h001C0011;14'd862:data <=32'h0016FFFA;14'd863:data <=32'h0009FFE6;
14'd864:data <=32'hFFF6FFD8;14'd865:data <=32'hFFE0FFD3;14'd866:data <=32'hFFCAFFD6;
14'd867:data <=32'hFFB7FFDE;14'd868:data <=32'hFFA9FFEB;14'd869:data <=32'hFFA0FFFB;
14'd870:data <=32'hFF9A0008;14'd871:data <=32'hFF960015;14'd872:data <=32'hFF930022;
14'd873:data <=32'hFF8F0030;14'd874:data <=32'hFF8A0041;14'd875:data <=32'hFF880056;
14'd876:data <=32'hFF8C0071;14'd877:data <=32'hFF97008D;14'd878:data <=32'hFFAB00A8;
14'd879:data <=32'hFFC900BD;14'd880:data <=32'hFFEC00CA;14'd881:data <=32'h001000CE;
14'd882:data <=32'h003400C7;14'd883:data <=32'h005300BA;14'd884:data <=32'h006E00A5;
14'd885:data <=32'h0082008D;14'd886:data <=32'h00900075;14'd887:data <=32'h0099005A;
14'd888:data <=32'h009C0040;14'd889:data <=32'h009A0027;14'd890:data <=32'h008F0010;
14'd891:data <=32'h0080FFFE;14'd892:data <=32'h006DFFF7;14'd893:data <=32'h005AFFF8;
14'd894:data <=32'h004E0004;14'd895:data <=32'h004C0014;14'd896:data <=32'h00E6002E;
14'd897:data <=32'h0100000A;14'd898:data <=32'h00F8FFDF;14'd899:data <=32'h007E0004;
14'd900:data <=32'h00A4003C;14'd901:data <=32'h00C00024;14'd902:data <=32'h00D50002;
14'd903:data <=32'h00E0FFD9;14'd904:data <=32'h00E0FFAF;14'd905:data <=32'h00D8FF85;
14'd906:data <=32'h00C6FF5C;14'd907:data <=32'h00ABFF37;14'd908:data <=32'h0087FF15;
14'd909:data <=32'h005AFEFC;14'd910:data <=32'h0026FEEF;14'd911:data <=32'hFFEFFEF1;
14'd912:data <=32'hFFBBFF01;14'd913:data <=32'hFF8FFF1F;14'd914:data <=32'hFF70FF46;
14'd915:data <=32'hFF5EFF70;14'd916:data <=32'hFF59FF98;14'd917:data <=32'hFF5DFFBA;
14'd918:data <=32'hFF66FFD5;14'd919:data <=32'hFF70FFEB;14'd920:data <=32'hFF7CFFFC;
14'd921:data <=32'hFF87000C;14'd922:data <=32'hFF94001A;14'd923:data <=32'hFFA40027;
14'd924:data <=32'hFFB70030;14'd925:data <=32'hFFCB0034;14'd926:data <=32'hFFDF0031;
14'd927:data <=32'hFFF20028;14'd928:data <=32'hFFFE001B;14'd929:data <=32'h0008000B;
14'd930:data <=32'h000BFFFA;14'd931:data <=32'h000AFFE9;14'd932:data <=32'h0005FFD9;
14'd933:data <=32'hFFFCFFCA;14'd934:data <=32'hFFEFFFBB;14'd935:data <=32'hFFDDFFAB;
14'd936:data <=32'hFFC4FFA0;14'd937:data <=32'hFFA5FF9D;14'd938:data <=32'hFF80FFA3;
14'd939:data <=32'hFF5BFFB5;14'd940:data <=32'hFF39FFD5;14'd941:data <=32'hFF220000;
14'd942:data <=32'hFF180033;14'd943:data <=32'hFF1E0068;14'd944:data <=32'hFF32009A;
14'd945:data <=32'hFF5400C4;14'd946:data <=32'hFF7D00E2;14'd947:data <=32'hFFAC00F4;
14'd948:data <=32'hFFDA00FA;14'd949:data <=32'h000700F6;14'd950:data <=32'h002F00E9;
14'd951:data <=32'h005300D5;14'd952:data <=32'h006F00BC;14'd953:data <=32'h0084009C;
14'd954:data <=32'h008F007B;14'd955:data <=32'h008F005A;14'd956:data <=32'h0086003F;
14'd957:data <=32'h0076002D;14'd958:data <=32'h00630026;14'd959:data <=32'h0055002A;
14'd960:data <=32'h003D0054;14'd961:data <=32'h004F0066;14'd962:data <=32'h006C005E;
14'd963:data <=32'h00910021;14'd964:data <=32'h00A90057;14'd965:data <=32'h00BA003E;
14'd966:data <=32'h00C50023;14'd967:data <=32'h00C70002;14'd968:data <=32'h00C3FFE6;
14'd969:data <=32'h00B9FFCC;14'd970:data <=32'h00ACFFB6;14'd971:data <=32'h009EFFA1;
14'd972:data <=32'h008EFF90;14'd973:data <=32'h007AFF81;14'd974:data <=32'h0063FF77;
14'd975:data <=32'h004BFF71;14'd976:data <=32'h0032FF71;14'd977:data <=32'h001EFF7A;
14'd978:data <=32'h000FFF86;14'd979:data <=32'h0007FF90;14'd980:data <=32'h0006FF99;
14'd981:data <=32'h0007FF9C;14'd982:data <=32'h0007FF99;14'd983:data <=32'h0001FF91;
14'd984:data <=32'hFFF5FF89;14'd985:data <=32'hFFE4FF86;14'd986:data <=32'hFFD0FF8A;
14'd987:data <=32'hFFBBFF94;14'd988:data <=32'hFFABFFA5;14'd989:data <=32'hFFA2FFBC;
14'd990:data <=32'hFFA0FFD2;14'd991:data <=32'hFFA5FFE7;14'd992:data <=32'hFFB0FFF8;
14'd993:data <=32'hFFBC0005;14'd994:data <=32'hFFCC000E;14'd995:data <=32'hFFDE0012;
14'd996:data <=32'hFFF20010;14'd997:data <=32'h00050007;14'd998:data <=32'h0014FFF7;
14'd999:data <=32'h001EFFE0;14'd1000:data <=32'h0021FFC4;14'd1001:data <=32'h0016FFA5;
14'd1002:data <=32'h0001FF89;14'd1003:data <=32'hFFDFFF75;14'd1004:data <=32'hFFB6FF6D;
14'd1005:data <=32'hFF8BFF73;14'd1006:data <=32'hFF64FF87;14'd1007:data <=32'hFF44FFA5;
14'd1008:data <=32'hFF2EFFCA;14'd1009:data <=32'hFF24FFF1;14'd1010:data <=32'hFF230018;
14'd1011:data <=32'hFF29003C;14'd1012:data <=32'hFF34005C;14'd1013:data <=32'hFF430079;
14'd1014:data <=32'hFF550092;14'd1015:data <=32'hFF6C00A9;14'd1016:data <=32'hFF8500BD;
14'd1017:data <=32'hFFA100CB;14'd1018:data <=32'hFFBF00D4;14'd1019:data <=32'hFFDB00D5;
14'd1020:data <=32'hFFF400D4;14'd1021:data <=32'h000900D2;14'd1022:data <=32'h001C00CF;
14'd1023:data <=32'h003100CF;14'd1024:data <=32'h002D0029;14'd1025:data <=32'h001B003A;
14'd1026:data <=32'h001F005D;14'd1027:data <=32'h007F00D7;14'd1028:data <=32'h00B60100;
14'd1029:data <=32'h00E300D6;14'd1030:data <=32'h010200A1;14'd1031:data <=32'h01140065;
14'd1032:data <=32'h0113002B;14'd1033:data <=32'h0103FFF8;14'd1034:data <=32'h00EBFFCC;
14'd1035:data <=32'h00CCFFAD;14'd1036:data <=32'h00AAFF96;14'd1037:data <=32'h0086FF88;
14'd1038:data <=32'h0063FF83;14'd1039:data <=32'h0042FF87;14'd1040:data <=32'h0024FF93;
14'd1041:data <=32'h000FFFA8;14'd1042:data <=32'h0004FFC3;14'd1043:data <=32'h0005FFDC;
14'd1044:data <=32'h0011FFF0;14'd1045:data <=32'h0024FFFB;14'd1046:data <=32'h003BFFFA;
14'd1047:data <=32'h004EFFEE;14'd1048:data <=32'h0059FFDA;14'd1049:data <=32'h005AFFC3;
14'd1050:data <=32'h0051FFAD;14'd1051:data <=32'h0043FF9C;14'd1052:data <=32'h002FFF92;
14'd1053:data <=32'h001CFF8F;14'd1054:data <=32'h0009FF90;14'd1055:data <=32'hFFFAFF96;
14'd1056:data <=32'hFFEDFF9D;14'd1057:data <=32'hFFE3FFA7;14'd1058:data <=32'hFFDBFFB2;
14'd1059:data <=32'hFFD7FFBF;14'd1060:data <=32'hFFD7FFCB;14'd1061:data <=32'hFFDBFFD7;
14'd1062:data <=32'hFFE4FFDF;14'd1063:data <=32'hFFF0FFE1;14'd1064:data <=32'hFFFCFFDD;
14'd1065:data <=32'h0005FFD2;14'd1066:data <=32'h0008FFC4;14'd1067:data <=32'h0004FFB4;
14'd1068:data <=32'hFFF9FFA7;14'd1069:data <=32'hFFEAFF9E;14'd1070:data <=32'hFFDBFF9B;
14'd1071:data <=32'hFFCCFF9D;14'd1072:data <=32'hFFBFFFA0;14'd1073:data <=32'hFFB6FFA5;
14'd1074:data <=32'hFFADFFA6;14'd1075:data <=32'hFFA4FFA4;14'd1076:data <=32'hFF95FFA3;
14'd1077:data <=32'hFF82FFA4;14'd1078:data <=32'hFF6AFFA8;14'd1079:data <=32'hFF4EFFB6;
14'd1080:data <=32'hFF36FFCA;14'd1081:data <=32'hFF20FFE7;14'd1082:data <=32'hFF100009;
14'd1083:data <=32'hFF050031;14'd1084:data <=32'hFF02005D;14'd1085:data <=32'hFF070089;
14'd1086:data <=32'hFF1300B8;14'd1087:data <=32'hFF2B00E9;14'd1088:data <=32'hFFED0071;
14'd1089:data <=32'hFFE0007C;14'd1090:data <=32'hFFC70093;14'd1091:data <=32'hFF76011A;
14'd1092:data <=32'hFFC00176;14'd1093:data <=32'h00100176;14'd1094:data <=32'h005B0160;
14'd1095:data <=32'h009B0139;14'd1096:data <=32'h00CA0104;14'd1097:data <=32'h00E900CC;
14'd1098:data <=32'h00F80092;14'd1099:data <=32'h00FB005E;14'd1100:data <=32'h00F3002C;
14'd1101:data <=32'h00E20000;14'd1102:data <=32'h00C9FFDC;14'd1103:data <=32'h00AAFFC0;
14'd1104:data <=32'h0087FFB0;14'd1105:data <=32'h0063FFAB;14'd1106:data <=32'h0044FFB0;
14'd1107:data <=32'h002CFFC0;14'd1108:data <=32'h0020FFD3;14'd1109:data <=32'h001CFFE5;
14'd1110:data <=32'h0022FFF3;14'd1111:data <=32'h002BFFFA;14'd1112:data <=32'h0034FFFA;
14'd1113:data <=32'h003BFFF6;14'd1114:data <=32'h003CFFEF;14'd1115:data <=32'h003BFFEA;
14'd1116:data <=32'h0038FFE8;14'd1117:data <=32'h0037FFE9;14'd1118:data <=32'h0038FFE8;
14'd1119:data <=32'h003DFFE8;14'd1120:data <=32'h0043FFE3;14'd1121:data <=32'h0047FFDC;
14'd1122:data <=32'h0049FFD2;14'd1123:data <=32'h0048FFC6;14'd1124:data <=32'h0044FFBC;
14'd1125:data <=32'h003DFFB2;14'd1126:data <=32'h0036FFAA;14'd1127:data <=32'h002EFFA3;
14'd1128:data <=32'h0026FF9D;14'd1129:data <=32'h001BFF97;14'd1130:data <=32'h000FFF91;
14'd1131:data <=32'hFFFFFF8E;14'd1132:data <=32'hFFF0FF91;14'd1133:data <=32'hFFDFFF99;
14'd1134:data <=32'hFFD3FFA5;14'd1135:data <=32'hFFCEFFB7;14'd1136:data <=32'hFFD1FFC5;
14'd1137:data <=32'hFFDBFFD1;14'd1138:data <=32'hFFEBFFD5;14'd1139:data <=32'hFFFBFFCE;
14'd1140:data <=32'h0008FFBC;14'd1141:data <=32'h000AFFA3;14'd1142:data <=32'h0000FF87;
14'd1143:data <=32'hFFECFF6E;14'd1144:data <=32'hFFCDFF5B;14'd1145:data <=32'hFFA6FF50;
14'd1146:data <=32'hFF7DFF4F;14'd1147:data <=32'hFF51FF5B;14'd1148:data <=32'hFF25FF70;
14'd1149:data <=32'hFEFDFF92;14'd1150:data <=32'hFEDAFFBE;14'd1151:data <=32'hFEBFFFF6;
14'd1152:data <=32'hFF3A000A;14'd1153:data <=32'hFF1A002E;14'd1154:data <=32'hFF070044;
14'd1155:data <=32'hFEE3003A;14'd1156:data <=32'hFEFD00B5;14'd1157:data <=32'hFF2900DD;
14'd1158:data <=32'hFF5C00F7;14'd1159:data <=32'hFF8F0105;14'd1160:data <=32'hFFBF0106;
14'd1161:data <=32'hFFE600FD;14'd1162:data <=32'h000800F2;14'd1163:data <=32'h002600E5;
14'd1164:data <=32'h004100D5;14'd1165:data <=32'h005A00C2;14'd1166:data <=32'h006F00AD;
14'd1167:data <=32'h00800093;14'd1168:data <=32'h008A0079;14'd1169:data <=32'h008F0060;
14'd1170:data <=32'h008E0048;14'd1171:data <=32'h008B0035;14'd1172:data <=32'h00880025;
14'd1173:data <=32'h00860016;14'd1174:data <=32'h00820006;14'd1175:data <=32'h007DFFF4;
14'd1176:data <=32'h0073FFE1;14'd1177:data <=32'h0064FFD0;14'd1178:data <=32'h004DFFC3;
14'd1179:data <=32'h0033FFC0;14'd1180:data <=32'h001AFFC6;14'd1181:data <=32'h0005FFD6;
14'd1182:data <=32'hFFF9FFEC;14'd1183:data <=32'hFFF70005;14'd1184:data <=32'hFFFF001C;
14'd1185:data <=32'h0010002E;14'd1186:data <=32'h00240037;14'd1187:data <=32'h003C0038;
14'd1188:data <=32'h00520033;14'd1189:data <=32'h00660028;14'd1190:data <=32'h00770017;
14'd1191:data <=32'h00840003;14'd1192:data <=32'h008BFFEB;14'd1193:data <=32'h008DFFD0;
14'd1194:data <=32'h0087FFB4;14'd1195:data <=32'h0079FF9A;14'd1196:data <=32'h0064FF84;
14'd1197:data <=32'h004AFF77;14'd1198:data <=32'h002EFF74;14'd1199:data <=32'h0015FF79;
14'd1200:data <=32'h0003FF86;14'd1201:data <=32'hFFF9FF96;14'd1202:data <=32'hFFFAFFA5;
14'd1203:data <=32'h0001FFAD;14'd1204:data <=32'h000BFFAC;14'd1205:data <=32'h0012FFA3;
14'd1206:data <=32'h0015FF94;14'd1207:data <=32'h000FFF81;14'd1208:data <=32'h0002FF70;
14'd1209:data <=32'hFFEEFF61;14'd1210:data <=32'hFFD6FF58;14'd1211:data <=32'hFFBBFF53;
14'd1212:data <=32'hFF9EFF53;14'd1213:data <=32'hFF7EFF59;14'd1214:data <=32'hFF5EFF66;
14'd1215:data <=32'hFF3EFF7B;14'd1216:data <=32'hFF7DFF1C;14'd1217:data <=32'hFF2FFF23;
14'd1218:data <=32'hFEFEFF48;14'd1219:data <=32'hFF44FFB0;14'd1220:data <=32'hFF460011;
14'd1221:data <=32'hFF550025;14'd1222:data <=32'hFF650031;14'd1223:data <=32'hFF750037;
14'd1224:data <=32'hFF7E0037;14'd1225:data <=32'hFF7F0038;14'd1226:data <=32'hFF7A003E;
14'd1227:data <=32'hFF75004A;14'd1228:data <=32'hFF72005F;14'd1229:data <=32'hFF750076;
14'd1230:data <=32'hFF810090;14'd1231:data <=32'hFF9400A7;14'd1232:data <=32'hFFAD00BA;
14'd1233:data <=32'hFFC900C8;14'd1234:data <=32'hFFE900D0;14'd1235:data <=32'h000B00D3;
14'd1236:data <=32'h002E00D0;14'd1237:data <=32'h005300C5;14'd1238:data <=32'h007600B0;
14'd1239:data <=32'h00940092;14'd1240:data <=32'h00A8006A;14'd1241:data <=32'h00B0003D;
14'd1242:data <=32'h00AA000F;14'd1243:data <=32'h0095FFE7;14'd1244:data <=32'h0076FFCB;
14'd1245:data <=32'h0051FFBD;14'd1246:data <=32'h002CFFBC;14'd1247:data <=32'h000CFFC8;
14'd1248:data <=32'hFFF6FFDC;14'd1249:data <=32'hFFE9FFF4;14'd1250:data <=32'hFFE4000C;
14'd1251:data <=32'hFFE70023;14'd1252:data <=32'hFFEF0038;14'd1253:data <=32'hFFFE0049;
14'd1254:data <=32'h000F0057;14'd1255:data <=32'h00260060;14'd1256:data <=32'h003F0063;
14'd1257:data <=32'h005A005F;14'd1258:data <=32'h00710053;14'd1259:data <=32'h00880042;
14'd1260:data <=32'h0096002B;14'd1261:data <=32'h00A00012;14'd1262:data <=32'h00A2FFFA;
14'd1263:data <=32'h00A0FFE4;14'd1264:data <=32'h009DFFD3;14'd1265:data <=32'h009BFFC3;
14'd1266:data <=32'h0099FFB2;14'd1267:data <=32'h0099FF9F;14'd1268:data <=32'h0096FF87;
14'd1269:data <=32'h008EFF6B;14'd1270:data <=32'h007DFF4D;14'd1271:data <=32'h0064FF33;
14'd1272:data <=32'h0040FF1C;14'd1273:data <=32'h0019FF11;14'd1274:data <=32'hFFF0FF0F;
14'd1275:data <=32'hFFC8FF18;14'd1276:data <=32'hFFA5FF28;14'd1277:data <=32'hFF87FF3C;
14'd1278:data <=32'hFF6EFF57;14'd1279:data <=32'hFF5CFF73;14'd1280:data <=32'h0047FF1F;
14'd1281:data <=32'h000BFEEE;14'd1282:data <=32'hFFBBFEE7;14'd1283:data <=32'hFF54FF99;
14'd1284:data <=32'hFF5FFFFC;14'd1285:data <=32'hFF7A0011;14'd1286:data <=32'hFF980017;
14'd1287:data <=32'hFFB30012;14'd1288:data <=32'hFFC40001;14'd1289:data <=32'hFFC7FFEB;
14'd1290:data <=32'hFFBFFFD7;14'd1291:data <=32'hFFABFFCC;14'd1292:data <=32'hFF91FFCC;
14'd1293:data <=32'hFF78FFD6;14'd1294:data <=32'hFF62FFE9;14'd1295:data <=32'hFF550003;
14'd1296:data <=32'hFF4E0022;14'd1297:data <=32'hFF4D0042;14'd1298:data <=32'hFF540062;
14'd1299:data <=32'hFF620082;14'd1300:data <=32'hFF7900A0;14'd1301:data <=32'hFF9800B8;
14'd1302:data <=32'hFFBE00C9;14'd1303:data <=32'hFFE900CF;14'd1304:data <=32'h001400C7;
14'd1305:data <=32'h003B00B3;14'd1306:data <=32'h00560095;14'd1307:data <=32'h00670073;
14'd1308:data <=32'h006C0051;14'd1309:data <=32'h00650033;14'd1310:data <=32'h0059001C;
14'd1311:data <=32'h004A000D;14'd1312:data <=32'h003B0003;14'd1313:data <=32'h002CFFFF;
14'd1314:data <=32'h001FFFFD;14'd1315:data <=32'h0013FFFB;14'd1316:data <=32'h0008FFFE;
14'd1317:data <=32'hFFFB0002;14'd1318:data <=32'hFFED000C;14'd1319:data <=32'hFFE3001A;
14'd1320:data <=32'hFFDE002D;14'd1321:data <=32'hFFDD0042;14'd1322:data <=32'hFFE40057;
14'd1323:data <=32'hFFF2006A;14'd1324:data <=32'h0003007B;14'd1325:data <=32'h00190089;
14'd1326:data <=32'h00320092;14'd1327:data <=32'h004F0098;14'd1328:data <=32'h0070009B;
14'd1329:data <=32'h00950095;14'd1330:data <=32'h00BC0088;14'd1331:data <=32'h00E5006E;
14'd1332:data <=32'h010A0047;14'd1333:data <=32'h01270013;14'd1334:data <=32'h0134FFD5;
14'd1335:data <=32'h0130FF92;14'd1336:data <=32'h011AFF52;14'd1337:data <=32'h00F2FF19;
14'd1338:data <=32'h00BEFEEE;14'd1339:data <=32'h0082FED3;14'd1340:data <=32'h0044FEC9;
14'd1341:data <=32'h0009FECB;14'd1342:data <=32'hFFD2FEDA;14'd1343:data <=32'hFFA3FEF3;
14'd1344:data <=32'h005CFF6E;14'd1345:data <=32'h0049FF41;14'd1346:data <=32'h001DFF10;
14'd1347:data <=32'hFF8BFF01;14'd1348:data <=32'hFF71FF6D;14'd1349:data <=32'hFF73FF92;
14'd1350:data <=32'hFF7DFFAF;14'd1351:data <=32'hFF8DFFC2;14'd1352:data <=32'hFF9DFFCA;
14'd1353:data <=32'hFFA7FFC8;14'd1354:data <=32'hFFAAFFC2;14'd1355:data <=32'hFFA4FFBE;
14'd1356:data <=32'hFF99FFBE;14'd1357:data <=32'hFF8DFFC5;14'd1358:data <=32'hFF82FFD1;
14'd1359:data <=32'hFF7BFFE0;14'd1360:data <=32'hFF77FFF1;14'd1361:data <=32'hFF78FFFF;
14'd1362:data <=32'hFF79000D;14'd1363:data <=32'hFF7B001D;14'd1364:data <=32'hFF81002C;
14'd1365:data <=32'hFF87003C;14'd1366:data <=32'hFF93004B;14'd1367:data <=32'hFFA10057;
14'd1368:data <=32'hFFB4005F;14'd1369:data <=32'hFFC60060;14'd1370:data <=32'hFFD6005C;
14'd1371:data <=32'hFFE10055;14'd1372:data <=32'hFFE6004E;14'd1373:data <=32'hFFE70049;
14'd1374:data <=32'hFFE80048;14'd1375:data <=32'hFFE9004C;14'd1376:data <=32'hFFEF0050;
14'd1377:data <=32'hFFFA0053;14'd1378:data <=32'h00070052;14'd1379:data <=32'h0015004B;
14'd1380:data <=32'h001D003E;14'd1381:data <=32'h0021002E;14'd1382:data <=32'h001E001E;
14'd1383:data <=32'h00140011;14'd1384:data <=32'h00050008;14'd1385:data <=32'hFFF30007;
14'd1386:data <=32'hFFE1000C;14'd1387:data <=32'hFFD00018;14'd1388:data <=32'hFFC40029;
14'd1389:data <=32'hFFBA0041;14'd1390:data <=32'hFFB8005B;14'd1391:data <=32'hFFBB007C;
14'd1392:data <=32'hFFCA009D;14'd1393:data <=32'hFFE200BE;14'd1394:data <=32'h000900DA;
14'd1395:data <=32'h003900EC;14'd1396:data <=32'h007300F0;14'd1397:data <=32'h00B000E1;
14'd1398:data <=32'h00E600C2;14'd1399:data <=32'h01150092;14'd1400:data <=32'h01330057;
14'd1401:data <=32'h01400018;14'd1402:data <=32'h013DFFDA;14'd1403:data <=32'h012CFFA2;
14'd1404:data <=32'h0110FF71;14'd1405:data <=32'h00EFFF49;14'd1406:data <=32'h00C9FF2B;
14'd1407:data <=32'h009FFF14;14'd1408:data <=32'h009AFF4B;14'd1409:data <=32'h0084FF26;
14'd1410:data <=32'h0074FF06;14'd1411:data <=32'h0094FEF9;14'd1412:data <=32'h0068FF34;
14'd1413:data <=32'h004EFF2E;14'd1414:data <=32'h0037FF29;14'd1415:data <=32'h0020FF27;
14'd1416:data <=32'h0009FF22;14'd1417:data <=32'hFFEDFF1D;14'd1418:data <=32'hFFCDFF1C;
14'd1419:data <=32'hFFA7FF22;14'd1420:data <=32'hFF82FF34;14'd1421:data <=32'hFF5EFF50;
14'd1422:data <=32'hFF46FF76;14'd1423:data <=32'hFF39FFA1;14'd1424:data <=32'hFF38FFCB;
14'd1425:data <=32'hFF42FFF2;14'd1426:data <=32'hFF550012;14'd1427:data <=32'hFF6A0029;
14'd1428:data <=32'hFF840038;14'd1429:data <=32'hFF9C0042;14'd1430:data <=32'hFFB40044;
14'd1431:data <=32'hFFCA0040;14'd1432:data <=32'hFFE00037;14'd1433:data <=32'hFFEF0029;
14'd1434:data <=32'hFFF70016;14'd1435:data <=32'hFFF70001;14'd1436:data <=32'hFFEDFFF0;
14'd1437:data <=32'hFFDCFFE4;14'd1438:data <=32'hFFC6FFE1;14'd1439:data <=32'hFFB2FFEA;
14'd1440:data <=32'hFFA3FFF9;14'd1441:data <=32'hFF9C000F;14'd1442:data <=32'hFF9E0025;
14'd1443:data <=32'hFFA80035;14'd1444:data <=32'hFFB60040;14'd1445:data <=32'hFFC60046;
14'd1446:data <=32'hFFD30044;14'd1447:data <=32'hFFDB003F;14'd1448:data <=32'hFFE0003A;
14'd1449:data <=32'hFFE00033;14'd1450:data <=32'hFFDC0030;14'd1451:data <=32'hFFD9002F;
14'd1452:data <=32'hFFD40030;14'd1453:data <=32'hFFCD0035;14'd1454:data <=32'hFFC5003C;
14'd1455:data <=32'hFFBF0047;14'd1456:data <=32'hFFBA0058;14'd1457:data <=32'hFFBA006E;
14'd1458:data <=32'hFFC10087;14'd1459:data <=32'hFFD200A1;14'd1460:data <=32'hFFEC00B6;
14'd1461:data <=32'h000F00C3;14'd1462:data <=32'h003300C6;14'd1463:data <=32'h005800BF;
14'd1464:data <=32'h007800AE;14'd1465:data <=32'h00900097;14'd1466:data <=32'h00A00081;
14'd1467:data <=32'h00AC006C;14'd1468:data <=32'h00B30058;14'd1469:data <=32'h00BD0047;
14'd1470:data <=32'h00C70036;14'd1471:data <=32'h00D10021;14'd1472:data <=32'h0129FFD3;
14'd1473:data <=32'h0129FF9A;14'd1474:data <=32'h0114FF7B;14'd1475:data <=32'h00F5FFFA;
14'd1476:data <=32'h00F6001E;14'd1477:data <=32'h0106FFF9;14'd1478:data <=32'h0110FFCE;
14'd1479:data <=32'h0111FF9D;14'd1480:data <=32'h0109FF69;14'd1481:data <=32'h00F1FF33;
14'd1482:data <=32'h00CBFF00;14'd1483:data <=32'h0096FED8;14'd1484:data <=32'h0053FEBD;
14'd1485:data <=32'h000CFEB7;14'd1486:data <=32'hFFC8FEC6;14'd1487:data <=32'hFF8CFEE7;
14'd1488:data <=32'hFF5EFF14;14'd1489:data <=32'hFF41FF48;14'd1490:data <=32'hFF33FF7E;
14'd1491:data <=32'hFF32FFB0;14'd1492:data <=32'hFF3BFFDD;14'd1493:data <=32'hFF4E0003;
14'd1494:data <=32'hFF680023;14'd1495:data <=32'hFF87003A;14'd1496:data <=32'hFFA90046;
14'd1497:data <=32'hFFCD0048;14'd1498:data <=32'hFFEC003E;14'd1499:data <=32'h0006002B;
14'd1500:data <=32'h00140011;14'd1501:data <=32'h0019FFF7;14'd1502:data <=32'h0011FFDE;
14'd1503:data <=32'h0002FFCC;14'd1504:data <=32'hFFF1FFC2;14'd1505:data <=32'hFFDEFFC0;
14'd1506:data <=32'hFFD0FFC2;14'd1507:data <=32'hFFC5FFC7;14'd1508:data <=32'hFFBCFFCC;
14'd1509:data <=32'hFFB3FFCF;14'd1510:data <=32'hFFA9FFD3;14'd1511:data <=32'hFF9FFFD6;
14'd1512:data <=32'hFF91FFDE;14'd1513:data <=32'hFF83FFEB;14'd1514:data <=32'hFF77FFFC;
14'd1515:data <=32'hFF700012;14'd1516:data <=32'hFF6E0029;14'd1517:data <=32'hFF71003F;
14'd1518:data <=32'hFF790054;14'd1519:data <=32'hFF840068;14'd1520:data <=32'hFF920079;
14'd1521:data <=32'hFFA10089;14'd1522:data <=32'hFFB30097;14'd1523:data <=32'hFFCA00A2;
14'd1524:data <=32'hFFE400A8;14'd1525:data <=32'hFFFE00A7;14'd1526:data <=32'h0018009F;
14'd1527:data <=32'h002E0090;14'd1528:data <=32'h003B007B;14'd1529:data <=32'h003E0066;
14'd1530:data <=32'h00380055;14'd1531:data <=32'h002B004D;14'd1532:data <=32'h001E0051;
14'd1533:data <=32'h0017005E;14'd1534:data <=32'h00190070;14'd1535:data <=32'h00250085;
14'd1536:data <=32'h00B600B3;14'd1537:data <=32'h00DF009B;14'd1538:data <=32'h00E70071;
14'd1539:data <=32'h00640074;14'd1540:data <=32'h007300B9;14'd1541:data <=32'h009B00B2;
14'd1542:data <=32'h00C700A0;14'd1543:data <=32'h00ED0083;14'd1544:data <=32'h01110059;
14'd1545:data <=32'h012A0023;14'd1546:data <=32'h0133FFE6;14'd1547:data <=32'h012BFFA5;
14'd1548:data <=32'h0110FF69;14'd1549:data <=32'h00E6FF38;14'd1550:data <=32'h00B2FF16;
14'd1551:data <=32'h007BFF06;14'd1552:data <=32'h0045FF04;14'd1553:data <=32'h0018FF0D;
14'd1554:data <=32'hFFEFFF1F;14'd1555:data <=32'hFFD0FF34;14'd1556:data <=32'hFFB6FF4C;
14'd1557:data <=32'hFFA1FF67;14'd1558:data <=32'hFF93FF84;14'd1559:data <=32'hFF8CFFA3;
14'd1560:data <=32'hFF8CFFC1;14'd1561:data <=32'hFF94FFDC;14'd1562:data <=32'hFFA2FFF2;
14'd1563:data <=32'hFFB50001;14'd1564:data <=32'hFFC70008;14'd1565:data <=32'hFFD7000A;
14'd1566:data <=32'hFFE60008;14'd1567:data <=32'hFFF10005;14'd1568:data <=32'hFFFC0001;
14'd1569:data <=32'h0004FFFC;14'd1570:data <=32'h000FFFF5;14'd1571:data <=32'h0019FFE9;
14'd1572:data <=32'h0022FFD8;14'd1573:data <=32'h0025FFC2;14'd1574:data <=32'h0020FFA7;
14'd1575:data <=32'h0011FF8C;14'd1576:data <=32'hFFF7FF76;14'd1577:data <=32'hFFD5FF67;
14'd1578:data <=32'hFFADFF64;14'd1579:data <=32'hFF85FF6D;14'd1580:data <=32'hFF60FF81;
14'd1581:data <=32'hFF41FF9F;14'd1582:data <=32'hFF2AFFC2;14'd1583:data <=32'hFF1DFFEB;
14'd1584:data <=32'hFF1A0014;14'd1585:data <=32'hFF1E003F;14'd1586:data <=32'hFF2D0068;
14'd1587:data <=32'hFF44008C;14'd1588:data <=32'hFF6500AA;14'd1589:data <=32'hFF8B00BD;
14'd1590:data <=32'hFFB600C5;14'd1591:data <=32'hFFDE00C0;14'd1592:data <=32'hFFFF00AF;
14'd1593:data <=32'h00150095;14'd1594:data <=32'h001E007B;14'd1595:data <=32'h001C0064;
14'd1596:data <=32'h00100056;14'd1597:data <=32'h00020053;14'd1598:data <=32'hFFF5005A;
14'd1599:data <=32'hFFF00069;14'd1600:data <=32'hFFE40087;14'd1601:data <=32'hFFF200A3;
14'd1602:data <=32'h001100A5;14'd1603:data <=32'h0039006E;14'd1604:data <=32'h003600B0;
14'd1605:data <=32'h004F00AE;14'd1606:data <=32'h006800A7;14'd1607:data <=32'h0082009D;
14'd1608:data <=32'h009C008C;14'd1609:data <=32'h00B30073;14'd1610:data <=32'h00C50054;
14'd1611:data <=32'h00CE002F;14'd1612:data <=32'h00CC000B;14'd1613:data <=32'h00C0FFEA;
14'd1614:data <=32'h00AEFFD2;14'd1615:data <=32'h0099FFC2;14'd1616:data <=32'h0086FFBA;
14'd1617:data <=32'h0078FFB7;14'd1618:data <=32'h006FFFB3;14'd1619:data <=32'h006AFFAF;
14'd1620:data <=32'h0064FFA5;14'd1621:data <=32'h005CFF9B;14'd1622:data <=32'h0050FF8F;
14'd1623:data <=32'h003FFF86;14'd1624:data <=32'h002DFF81;14'd1625:data <=32'h0019FF80;
14'd1626:data <=32'h0008FF85;14'd1627:data <=32'hFFF7FF8A;14'd1628:data <=32'hFFE8FF93;
14'd1629:data <=32'hFFDAFF9E;14'd1630:data <=32'hFFCEFFAD;14'd1631:data <=32'hFFC5FFBE;
14'd1632:data <=32'hFFC1FFD4;14'd1633:data <=32'hFFC4FFEB;14'd1634:data <=32'hFFD10001;
14'd1635:data <=32'hFFE70012;14'd1636:data <=32'h0003001A;14'd1637:data <=32'h00210015;
14'd1638:data <=32'h003C0003;14'd1639:data <=32'h0051FFE7;14'd1640:data <=32'h0059FFC3;
14'd1641:data <=32'h0054FF9D;14'd1642:data <=32'h0043FF7B;14'd1643:data <=32'h0028FF61;
14'd1644:data <=32'h0006FF4D;14'd1645:data <=32'hFFE0FF44;14'd1646:data <=32'hFFBAFF45;
14'd1647:data <=32'hFF95FF4C;14'd1648:data <=32'hFF73FF5C;14'd1649:data <=32'hFF54FF74;
14'd1650:data <=32'hFF3AFF90;14'd1651:data <=32'hFF26FFB4;14'd1652:data <=32'hFF1DFFDB;
14'd1653:data <=32'hFF1C0002;14'd1654:data <=32'hFF250026;14'd1655:data <=32'hFF350043;
14'd1656:data <=32'hFF4A005A;14'd1657:data <=32'hFF5C0066;14'd1658:data <=32'hFF6C0070;
14'd1659:data <=32'hFF760077;14'd1660:data <=32'hFF7E0081;14'd1661:data <=32'hFF83008F;
14'd1662:data <=32'hFF8D00A2;14'd1663:data <=32'hFF9D00B6;14'd1664:data <=32'hFFDE001F;
14'd1665:data <=32'hFFC5002D;14'd1666:data <=32'hFFBB0050;14'd1667:data <=32'hFFF100D9;
14'd1668:data <=32'h00070116;14'd1669:data <=32'h00370108;14'd1670:data <=32'h006000F2;
14'd1671:data <=32'h008000D4;14'd1672:data <=32'h009B00B3;14'd1673:data <=32'h00AF008E;
14'd1674:data <=32'h00B90064;14'd1675:data <=32'h00B7003C;14'd1676:data <=32'h00AA0015;
14'd1677:data <=32'h0092FFF8;14'd1678:data <=32'h0074FFE6;14'd1679:data <=32'h0056FFE1;
14'd1680:data <=32'h003DFFE9;14'd1681:data <=32'h002DFFFA;14'd1682:data <=32'h002A000F;
14'd1683:data <=32'h0031001E;14'd1684:data <=32'h00400028;14'd1685:data <=32'h00520029;
14'd1686:data <=32'h00630021;14'd1687:data <=32'h00700012;14'd1688:data <=32'h00780001;
14'd1689:data <=32'h007DFFEE;14'd1690:data <=32'h007BFFDB;14'd1691:data <=32'h0076FFC8;
14'd1692:data <=32'h006CFFB4;14'd1693:data <=32'h005CFFA4;14'd1694:data <=32'h0047FF97;
14'd1695:data <=32'h002FFF92;14'd1696:data <=32'h0017FF93;14'd1697:data <=32'h0000FF9F;
14'd1698:data <=32'hFFF0FFB1;14'd1699:data <=32'hFFE9FFC7;14'd1700:data <=32'hFFEBFFDD;
14'd1701:data <=32'hFFF7FFEE;14'd1702:data <=32'h0009FFF7;14'd1703:data <=32'h001BFFF9;
14'd1704:data <=32'h002DFFF2;14'd1705:data <=32'h0038FFE4;14'd1706:data <=32'h003EFFD4;
14'd1707:data <=32'h003FFFC4;14'd1708:data <=32'h003CFFB5;14'd1709:data <=32'h0038FFA9;
14'd1710:data <=32'h0032FF9C;14'd1711:data <=32'h002DFF8F;14'd1712:data <=32'h0023FF81;
14'd1713:data <=32'h0016FF72;14'd1714:data <=32'h0006FF65;14'd1715:data <=32'hFFF1FF59;
14'd1716:data <=32'hFFD7FF52;14'd1717:data <=32'hFFBDFF4F;14'd1718:data <=32'hFFA1FF50;
14'd1719:data <=32'hFF87FF56;14'd1720:data <=32'hFF6CFF5E;14'd1721:data <=32'hFF4FFF69;
14'd1722:data <=32'hFF2FFF79;14'd1723:data <=32'hFF0EFF91;14'd1724:data <=32'hFEEDFFB2;
14'd1725:data <=32'hFED1FFE1;14'd1726:data <=32'hFEC0001A;14'd1727:data <=32'hFEBF005A;
14'd1728:data <=32'hFFB8002F;14'd1729:data <=32'hFFA5002F;14'd1730:data <=32'hFF7F0038;
14'd1731:data <=32'hFF0000A6;14'd1732:data <=32'hFF1A0111;14'd1733:data <=32'hFF580130;
14'd1734:data <=32'hFF99013D;14'd1735:data <=32'hFFD8013C;14'd1736:data <=32'h0014012E;
14'd1737:data <=32'h00490115;14'd1738:data <=32'h007500EF;14'd1739:data <=32'h009600C1;
14'd1740:data <=32'h00A6008F;14'd1741:data <=32'h00A6005D;14'd1742:data <=32'h00980033;
14'd1743:data <=32'h007F0014;14'd1744:data <=32'h00620003;14'd1745:data <=32'h00470000;
14'd1746:data <=32'h00330006;14'd1747:data <=32'h00270013;14'd1748:data <=32'h0025001E;
14'd1749:data <=32'h00270027;14'd1750:data <=32'h002D002A;14'd1751:data <=32'h0034002C;
14'd1752:data <=32'h0039002C;14'd1753:data <=32'h003E0029;14'd1754:data <=32'h00440028;
14'd1755:data <=32'h004A0024;14'd1756:data <=32'h0052001F;14'd1757:data <=32'h00580017;
14'd1758:data <=32'h005C000C;14'd1759:data <=32'h005C0000;14'd1760:data <=32'h0059FFF6;
14'd1761:data <=32'h0054FFEE;14'd1762:data <=32'h004EFFE9;14'd1763:data <=32'h0049FFE7;
14'd1764:data <=32'h0048FFE7;14'd1765:data <=32'h004AFFE6;14'd1766:data <=32'h004CFFE1;
14'd1767:data <=32'h004FFFD9;14'd1768:data <=32'h004DFFCD;14'd1769:data <=32'h0047FFC1;
14'd1770:data <=32'h003CFFB8;14'd1771:data <=32'h002FFFB5;14'd1772:data <=32'h0021FFB8;
14'd1773:data <=32'h0018FFC0;14'd1774:data <=32'h0014FFCC;14'd1775:data <=32'h0018FFD8;
14'd1776:data <=32'h0023FFDE;14'd1777:data <=32'h0033FFE0;14'd1778:data <=32'h0043FFD8;
14'd1779:data <=32'h0051FFCA;14'd1780:data <=32'h005CFFB5;14'd1781:data <=32'h0060FF9A;
14'd1782:data <=32'h005FFF7D;14'd1783:data <=32'h0056FF5D;14'd1784:data <=32'h0045FF3A;
14'd1785:data <=32'h0029FF19;14'd1786:data <=32'h0000FEFB;14'd1787:data <=32'hFFCCFEE7;
14'd1788:data <=32'hFF8DFEDF;14'd1789:data <=32'hFF48FEEB;14'd1790:data <=32'hFF06FF0A;
14'd1791:data <=32'hFECEFF3E;14'd1792:data <=32'hFF55FF9F;14'd1793:data <=32'hFF30FFAE;
14'd1794:data <=32'hFF15FFB0;14'd1795:data <=32'hFEE1FF91;14'd1796:data <=32'hFEC30007;
14'd1797:data <=32'hFED2003C;14'd1798:data <=32'hFEEA006B;14'd1799:data <=32'hFF080090;
14'd1800:data <=32'hFF2A00B1;14'd1801:data <=32'hFF5200C9;14'd1802:data <=32'hFF7D00D8;
14'd1803:data <=32'hFFA700DC;14'd1804:data <=32'hFFCE00D5;14'd1805:data <=32'hFFEE00C8;
14'd1806:data <=32'h000600B6;14'd1807:data <=32'h001500A5;14'd1808:data <=32'h00200095;
14'd1809:data <=32'h0028008C;14'd1810:data <=32'h00310084;14'd1811:data <=32'h003D007D;
14'd1812:data <=32'h004B0071;14'd1813:data <=32'h00590062;14'd1814:data <=32'h0062004D;
14'd1815:data <=32'h00630036;14'd1816:data <=32'h005E001F;14'd1817:data <=32'h0052000D;
14'd1818:data <=32'h00420001;14'd1819:data <=32'h0030FFFC;14'd1820:data <=32'h0020FFFF;
14'd1821:data <=32'h00130005;14'd1822:data <=32'h000B000F;14'd1823:data <=32'h0006001A;
14'd1824:data <=32'h00040026;14'd1825:data <=32'h00070033;14'd1826:data <=32'h000E0041;
14'd1827:data <=32'h001A004D;14'd1828:data <=32'h002C0056;14'd1829:data <=32'h0043005A;
14'd1830:data <=32'h005D0055;14'd1831:data <=32'h00740047;14'd1832:data <=32'h0087002F;
14'd1833:data <=32'h00910013;14'd1834:data <=32'h0090FFF6;14'd1835:data <=32'h0086FFDC;
14'd1836:data <=32'h0075FFCA;14'd1837:data <=32'h0060FFC0;14'd1838:data <=32'h004DFFBF;
14'd1839:data <=32'h003FFFC6;14'd1840:data <=32'h0039FFCF;14'd1841:data <=32'h003AFFD8;
14'd1842:data <=32'h003FFFDE;14'd1843:data <=32'h0049FFE0;14'd1844:data <=32'h0055FFDD;
14'd1845:data <=32'h0060FFD3;14'd1846:data <=32'h006BFFC6;14'd1847:data <=32'h0075FFB3;
14'd1848:data <=32'h007AFF9B;14'd1849:data <=32'h007BFF7D;14'd1850:data <=32'h0072FF59;
14'd1851:data <=32'h005DFF36;14'd1852:data <=32'h003EFF16;14'd1853:data <=32'h0011FEFE;
14'd1854:data <=32'hFFDDFEF3;14'd1855:data <=32'hFFA7FEFA;14'd1856:data <=32'hFFF6FEE5;
14'd1857:data <=32'hFFB1FECE;14'd1858:data <=32'hFF80FED5;14'd1859:data <=32'hFFA0FF34;
14'd1860:data <=32'hFF75FF84;14'd1861:data <=32'hFF70FF93;14'd1862:data <=32'hFF6BFFA0;
14'd1863:data <=32'hFF64FFAA;14'd1864:data <=32'hFF58FFB7;14'd1865:data <=32'hFF4FFFC8;
14'd1866:data <=32'hFF45FFDB;14'd1867:data <=32'hFF40FFF1;14'd1868:data <=32'hFF3D0006;
14'd1869:data <=32'hFF3D001E;14'd1870:data <=32'hFF3C0035;14'd1871:data <=32'hFF3E0050;
14'd1872:data <=32'hFF45006D;14'd1873:data <=32'hFF53008E;14'd1874:data <=32'hFF6A00AE;
14'd1875:data <=32'hFF8D00CA;14'd1876:data <=32'hFFB900DC;14'd1877:data <=32'hFFE900E1;
14'd1878:data <=32'h001900D6;14'd1879:data <=32'h004300BD;14'd1880:data <=32'h0062009A;
14'd1881:data <=32'h00720074;14'd1882:data <=32'h0076004B;14'd1883:data <=32'h006F0027;
14'd1884:data <=32'h005F000B;14'd1885:data <=32'h004AFFF6;14'd1886:data <=32'h0032FFE8;
14'd1887:data <=32'h0018FFE3;14'd1888:data <=32'hFFFFFFE6;14'd1889:data <=32'hFFE8FFEF;
14'd1890:data <=32'hFFD30001;14'd1891:data <=32'hFFC7001A;14'd1892:data <=32'hFFC30035;
14'd1893:data <=32'hFFCA0052;14'd1894:data <=32'hFFDA006B;14'd1895:data <=32'hFFF3007D;
14'd1896:data <=32'h000F0087;14'd1897:data <=32'h002B0087;14'd1898:data <=32'h0044007E;
14'd1899:data <=32'h00570071;14'd1900:data <=32'h00650063;14'd1901:data <=32'h006D0056;
14'd1902:data <=32'h0075004C;14'd1903:data <=32'h007E0044;14'd1904:data <=32'h0089003D;
14'd1905:data <=32'h00960032;14'd1906:data <=32'h00A40022;14'd1907:data <=32'h00AF000D;
14'd1908:data <=32'h00B7FFF5;14'd1909:data <=32'h00B8FFDA;14'd1910:data <=32'h00B6FFBF;
14'd1911:data <=32'h00AFFFA6;14'd1912:data <=32'h00A4FF8D;14'd1913:data <=32'h0095FF76;
14'd1914:data <=32'h0084FF60;14'd1915:data <=32'h006EFF4B;14'd1916:data <=32'h0052FF3A;
14'd1917:data <=32'h0030FF2F;14'd1918:data <=32'h000CFF2D;14'd1919:data <=32'hFFE9FF34;
14'd1920:data <=32'h00C7FF47;14'd1921:data <=32'h00A8FF03;14'd1922:data <=32'h006AFEDF;
14'd1923:data <=32'hFFDDFF61;14'd1924:data <=32'hFFC2FFB0;14'd1925:data <=32'hFFD2FFBB;
14'd1926:data <=32'hFFE2FFBA;14'd1927:data <=32'hFFEFFFAF;14'd1928:data <=32'hFFF1FF9F;
14'd1929:data <=32'hFFEBFF90;14'd1930:data <=32'hFFDDFF80;14'd1931:data <=32'hFFCAFF76;
14'd1932:data <=32'hFFB3FF70;14'd1933:data <=32'hFF97FF70;14'd1934:data <=32'hFF78FF75;
14'd1935:data <=32'hFF56FF84;14'd1936:data <=32'hFF37FF9D;14'd1937:data <=32'hFF1DFFC2;
14'd1938:data <=32'hFF0CFFF1;14'd1939:data <=32'hFF0B0024;14'd1940:data <=32'hFF1A0058;
14'd1941:data <=32'hFF380084;14'd1942:data <=32'hFF6000A3;14'd1943:data <=32'hFF8D00B5;
14'd1944:data <=32'hFFBA00B9;14'd1945:data <=32'hFFE300AF;14'd1946:data <=32'h0002009F;
14'd1947:data <=32'h001A008A;14'd1948:data <=32'h002C0072;14'd1949:data <=32'h00360059;
14'd1950:data <=32'h003B0043;14'd1951:data <=32'h003A002B;14'd1952:data <=32'h00330014;
14'd1953:data <=32'h00270002;14'd1954:data <=32'h0016FFF4;14'd1955:data <=32'h0000FFED;
14'd1956:data <=32'hFFEAFFEE;14'd1957:data <=32'hFFD6FFF6;14'd1958:data <=32'hFFC60004;
14'd1959:data <=32'hFFBB0015;14'd1960:data <=32'hFFB60026;14'd1961:data <=32'hFFB40038;
14'd1962:data <=32'hFFB4004A;14'd1963:data <=32'hFFB6005C;14'd1964:data <=32'hFFB90070;
14'd1965:data <=32'hFFC00089;14'd1966:data <=32'hFFCF00A3;14'd1967:data <=32'hFFE600BE;
14'd1968:data <=32'h000800D5;14'd1969:data <=32'h003300E5;14'd1970:data <=32'h006600E8;
14'd1971:data <=32'h009900DC;14'd1972:data <=32'h00CC00C3;14'd1973:data <=32'h00F5009C;
14'd1974:data <=32'h0113006D;14'd1975:data <=32'h01260038;14'd1976:data <=32'h012C0001;
14'd1977:data <=32'h0127FFCA;14'd1978:data <=32'h0117FF95;14'd1979:data <=32'h00FBFF66;
14'd1980:data <=32'h00D5FF3D;14'd1981:data <=32'h00A6FF1D;14'd1982:data <=32'h0071FF0D;
14'd1983:data <=32'h003BFF0C;14'd1984:data <=32'h00B3FFCA;14'd1985:data <=32'h00BCFF9C;
14'd1986:data <=32'h00AFFF61;14'd1987:data <=32'h0026FF22;14'd1988:data <=32'hFFF2FF74;
14'd1989:data <=32'hFFF1FF89;14'd1990:data <=32'hFFF7FF97;14'd1991:data <=32'hFFFFFF9B;
14'd1992:data <=32'h0004FF99;14'd1993:data <=32'h0005FF95;14'd1994:data <=32'h0000FF8E;
14'd1995:data <=32'hFFF9FF87;14'd1996:data <=32'hFFF0FF81;14'd1997:data <=32'hFFE4FF7B;
14'd1998:data <=32'hFFD5FF76;14'd1999:data <=32'hFFC1FF73;14'd2000:data <=32'hFFA9FF75;
14'd2001:data <=32'hFF8FFF7F;14'd2002:data <=32'hFF78FF91;14'd2003:data <=32'hFF65FFAC;
14'd2004:data <=32'hFF5BFFCA;14'd2005:data <=32'hFF5DFFE9;14'd2006:data <=32'hFF660005;
14'd2007:data <=32'hFF750019;14'd2008:data <=32'hFF860026;14'd2009:data <=32'hFF95002C;
14'd2010:data <=32'hFFA00030;14'd2011:data <=32'hFFA70033;14'd2012:data <=32'hFFAE0037;
14'd2013:data <=32'hFFB6003E;14'd2014:data <=32'hFFC00043;14'd2015:data <=32'hFFCD0048;
14'd2016:data <=32'hFFDB0049;14'd2017:data <=32'hFFE80044;14'd2018:data <=32'hFFF5003C;
14'd2019:data <=32'hFFFD0032;14'd2020:data <=32'h00020025;14'd2021:data <=32'h00010019;
14'd2022:data <=32'hFFFE000D;14'd2023:data <=32'hFFF90002;14'd2024:data <=32'hFFEFFFF7;
14'd2025:data <=32'hFFE1FFEE;14'd2026:data <=32'hFFCFFFE8;14'd2027:data <=32'hFFB6FFE8;
14'd2028:data <=32'hFF9AFFF0;14'd2029:data <=32'hFF7E0004;14'd2030:data <=32'hFF660024;
14'd2031:data <=32'hFF58004F;14'd2032:data <=32'hFF580081;14'd2033:data <=32'hFF6700B5;
14'd2034:data <=32'hFF8800E5;14'd2035:data <=32'hFFB60109;14'd2036:data <=32'hFFEF0120;
14'd2037:data <=32'h002B0128;14'd2038:data <=32'h00680120;14'd2039:data <=32'h009E010B;
14'd2040:data <=32'h00D000EA;14'd2041:data <=32'h00F800C0;14'd2042:data <=32'h01170091;
14'd2043:data <=32'h012A005A;14'd2044:data <=32'h01310021;14'd2045:data <=32'h0129FFE9;
14'd2046:data <=32'h0115FFB4;14'd2047:data <=32'h00F4FF8B;14'd2048:data <=32'h00C3FFC9;
14'd2049:data <=32'h00C2FFAC;14'd2050:data <=32'h00C8FF92;14'd2051:data <=32'h00F2FF82;
14'd2052:data <=32'h00BEFFA9;14'd2053:data <=32'h00B7FF98;14'd2054:data <=32'h00ADFF84;
14'd2055:data <=32'h00A3FF6C;14'd2056:data <=32'h008EFF52;14'd2057:data <=32'h0073FF3E;
14'd2058:data <=32'h0051FF30;14'd2059:data <=32'h002DFF29;14'd2060:data <=32'h000AFF2C;
14'd2061:data <=32'hFFEAFF35;14'd2062:data <=32'hFFCEFF44;14'd2063:data <=32'hFFB7FF56;
14'd2064:data <=32'hFFA3FF6A;14'd2065:data <=32'hFF94FF82;14'd2066:data <=32'hFF89FF9C;
14'd2067:data <=32'hFF85FFBA;14'd2068:data <=32'hFF8AFFD7;14'd2069:data <=32'hFF97FFEF;
14'd2070:data <=32'hFFAC0000;14'd2071:data <=32'hFFC30007;14'd2072:data <=32'hFFD90002;
14'd2073:data <=32'hFFE8FFF7;14'd2074:data <=32'hFFEDFFE4;14'd2075:data <=32'hFFE9FFD5;
14'd2076:data <=32'hFFDEFFC9;14'd2077:data <=32'hFFCEFFC5;14'd2078:data <=32'hFFBDFFC9;
14'd2079:data <=32'hFFB1FFD2;14'd2080:data <=32'hFFA8FFDF;14'd2081:data <=32'hFFA5FFED;
14'd2082:data <=32'hFFA6FFFA;14'd2083:data <=32'hFFAA0006;14'd2084:data <=32'hFFB0000F;
14'd2085:data <=32'hFFB70016;14'd2086:data <=32'hFFC1001B;14'd2087:data <=32'hFFCC001C;
14'd2088:data <=32'hFFD40019;14'd2089:data <=32'hFFDC0010;14'd2090:data <=32'hFFDE0004;
14'd2091:data <=32'hFFD9FFF6;14'd2092:data <=32'hFFCCFFE9;14'd2093:data <=32'hFFB7FFE2;
14'd2094:data <=32'hFF9DFFE4;14'd2095:data <=32'hFF82FFF1;14'd2096:data <=32'hFF6C000A;
14'd2097:data <=32'hFF5E002B;14'd2098:data <=32'hFF5B0050;14'd2099:data <=32'hFF640076;
14'd2100:data <=32'hFF760096;14'd2101:data <=32'hFF8E00AF;14'd2102:data <=32'hFFAB00C4;
14'd2103:data <=32'hFFC800D1;14'd2104:data <=32'hFFE500DA;14'd2105:data <=32'h000300DE;
14'd2106:data <=32'h002200DF;14'd2107:data <=32'h004300DC;14'd2108:data <=32'h006200D2;
14'd2109:data <=32'h007F00C4;14'd2110:data <=32'h009800AF;14'd2111:data <=32'h00AC0099;
14'd2112:data <=32'h00FF005A;14'd2113:data <=32'h010B0031;14'd2114:data <=32'h0103001E;
14'd2115:data <=32'h00D00095;14'd2116:data <=32'h00CB00BB;14'd2117:data <=32'h00F7009F;
14'd2118:data <=32'h011D0078;14'd2119:data <=32'h013C0042;14'd2120:data <=32'h014C0002;
14'd2121:data <=32'h0147FFBE;14'd2122:data <=32'h0131FF7F;14'd2123:data <=32'h010CFF47;
14'd2124:data <=32'h00DAFF1D;14'd2125:data <=32'h00A5FF01;14'd2126:data <=32'h006BFEF4;
14'd2127:data <=32'h0034FEF3;14'd2128:data <=32'hFFFFFEFD;14'd2129:data <=32'hFFCEFF13;
14'd2130:data <=32'hFFA7FF33;14'd2131:data <=32'hFF89FF5D;14'd2132:data <=32'hFF78FF8A;
14'd2133:data <=32'hFF77FFBA;14'd2134:data <=32'hFF85FFE3;14'd2135:data <=32'hFF9E0003;
14'd2136:data <=32'hFFBF0015;14'd2137:data <=32'hFFDE001A;14'd2138:data <=32'hFFFB0013;
14'd2139:data <=32'h000D0003;14'd2140:data <=32'h0018FFF0;14'd2141:data <=32'h001AFFDE;
14'd2142:data <=32'h0016FFCF;14'd2143:data <=32'h000FFFC3;14'd2144:data <=32'h0007FFBA;
14'd2145:data <=32'hFFFEFFB4;14'd2146:data <=32'hFFF5FFAF;14'd2147:data <=32'hFFEBFFAB;
14'd2148:data <=32'hFFDFFFA8;14'd2149:data <=32'hFFD1FFA8;14'd2150:data <=32'hFFC4FFAB;
14'd2151:data <=32'hFFB7FFB0;14'd2152:data <=32'hFFADFFB9;14'd2153:data <=32'hFFA6FFC0;
14'd2154:data <=32'hFF9FFFC8;14'd2155:data <=32'hFF99FFCE;14'd2156:data <=32'hFF92FFD5;
14'd2157:data <=32'hFF88FFDB;14'd2158:data <=32'hFF7EFFE6;14'd2159:data <=32'hFF73FFF5;
14'd2160:data <=32'hFF6C000B;14'd2161:data <=32'hFF6B0022;14'd2162:data <=32'hFF72003B;
14'd2163:data <=32'hFF7F004F;14'd2164:data <=32'hFF92005D;14'd2165:data <=32'hFFA50062;
14'd2166:data <=32'hFFB50061;14'd2167:data <=32'hFFC0005D;14'd2168:data <=32'hFFC40056;
14'd2169:data <=32'hFFC10053;14'd2170:data <=32'hFFBB0056;14'd2171:data <=32'hFFB5005E;
14'd2172:data <=32'hFFB1006B;14'd2173:data <=32'hFFB2007D;14'd2174:data <=32'hFFB60091;
14'd2175:data <=32'hFFBD00A6;14'd2176:data <=32'h004300EC;14'd2177:data <=32'h006700E9;
14'd2178:data <=32'h007000D1;14'd2179:data <=32'hFFEB00C0;14'd2180:data <=32'hFFE60112;
14'd2181:data <=32'h001F0126;14'd2182:data <=32'h005F012A;14'd2183:data <=32'h00A1011C;
14'd2184:data <=32'h00DD00F9;14'd2185:data <=32'h010D00C6;14'd2186:data <=32'h012D0089;
14'd2187:data <=32'h013B0049;14'd2188:data <=32'h0138000B;14'd2189:data <=32'h012BFFD3;
14'd2190:data <=32'h0112FFA1;14'd2191:data <=32'h00F0FF78;14'd2192:data <=32'h00CBFF57;
14'd2193:data <=32'h009EFF40;14'd2194:data <=32'h006EFF34;14'd2195:data <=32'h0040FF34;
14'd2196:data <=32'h0015FF40;14'd2197:data <=32'hFFF1FF56;14'd2198:data <=32'hFFD9FF73;
14'd2199:data <=32'hFFCDFF92;14'd2200:data <=32'hFFC9FFAF;14'd2201:data <=32'hFFCEFFC5;
14'd2202:data <=32'hFFD6FFD4;14'd2203:data <=32'hFFDEFFDF;14'd2204:data <=32'hFFE5FFE6;
14'd2205:data <=32'hFFEBFFEE;14'd2206:data <=32'hFFF1FFF4;14'd2207:data <=32'hFFFBFFFB;
14'd2208:data <=32'h00080001;14'd2209:data <=32'h00190001;14'd2210:data <=32'h002AFFFC;
14'd2211:data <=32'h003BFFEF;14'd2212:data <=32'h0047FFDB;14'd2213:data <=32'h004DFFC4;
14'd2214:data <=32'h004AFFAA;14'd2215:data <=32'h0040FF8F;14'd2216:data <=32'h002FFF7A;
14'd2217:data <=32'h0019FF68;14'd2218:data <=32'hFFFFFF59;14'd2219:data <=32'hFFE1FF51;
14'd2220:data <=32'hFFC0FF4E;14'd2221:data <=32'hFF9EFF53;14'd2222:data <=32'hFF7AFF60;
14'd2223:data <=32'hFF59FF78;14'd2224:data <=32'hFF3EFF9A;14'd2225:data <=32'hFF2EFFC3;
14'd2226:data <=32'hFF2AFFEF;14'd2227:data <=32'hFF340018;14'd2228:data <=32'hFF4B003B;
14'd2229:data <=32'hFF680051;14'd2230:data <=32'hFF87005B;14'd2231:data <=32'hFFA2005A;
14'd2232:data <=32'hFFB5004F;14'd2233:data <=32'hFFC00042;14'd2234:data <=32'hFFC20035;
14'd2235:data <=32'hFFBC002C;14'd2236:data <=32'hFFB30028;14'd2237:data <=32'hFFA60028;
14'd2238:data <=32'hFF990030;14'd2239:data <=32'hFF8C003F;14'd2240:data <=32'hFF8A005F;
14'd2241:data <=32'hFF80007C;14'd2242:data <=32'hFF8E008B;14'd2243:data <=32'hFFB00064;
14'd2244:data <=32'hFF8F00B4;14'd2245:data <=32'hFFA900D0;14'd2246:data <=32'hFFCF00E6;
14'd2247:data <=32'hFFF900F1;14'd2248:data <=32'h002600EF;14'd2249:data <=32'h004F00DF;
14'd2250:data <=32'h007000C7;14'd2251:data <=32'h008800AB;14'd2252:data <=32'h0097008E;
14'd2253:data <=32'h00A00075;14'd2254:data <=32'h00A5005D;14'd2255:data <=32'h00A80047;
14'd2256:data <=32'h00AB0032;14'd2257:data <=32'h00AB001C;14'd2258:data <=32'h00A70006;
14'd2259:data <=32'h00A1FFF1;14'd2260:data <=32'h0095FFDE;14'd2261:data <=32'h0089FFCF;
14'd2262:data <=32'h007CFFC5;14'd2263:data <=32'h0072FFBC;14'd2264:data <=32'h0067FFB4;
14'd2265:data <=32'h005CFFAA;14'd2266:data <=32'h004EFFA0;14'd2267:data <=32'h003CFF97;
14'd2268:data <=32'h0026FF93;14'd2269:data <=32'h000CFF96;14'd2270:data <=32'hFFF5FFA3;
14'd2271:data <=32'hFFE0FFB7;14'd2272:data <=32'hFFD7FFD2;14'd2273:data <=32'hFFD8FFF0;
14'd2274:data <=32'hFFE4000A;14'd2275:data <=32'hFFFB001D;14'd2276:data <=32'h00170027;
14'd2277:data <=32'h00340026;14'd2278:data <=32'h0050001B;14'd2279:data <=32'h00660007;
14'd2280:data <=32'h0077FFEE;14'd2281:data <=32'h0082FFD0;14'd2282:data <=32'h0084FFAE;
14'd2283:data <=32'h007DFF8B;14'd2284:data <=32'h006EFF69;14'd2285:data <=32'h0054FF4A;
14'd2286:data <=32'h0032FF32;14'd2287:data <=32'h0008FF23;14'd2288:data <=32'hFFDCFF1F;
14'd2289:data <=32'hFFB0FF2A;14'd2290:data <=32'hFF89FF3F;14'd2291:data <=32'hFF6EFF5E;
14'd2292:data <=32'hFF5CFF7E;14'd2293:data <=32'hFF56FF9D;14'd2294:data <=32'hFF57FFB6;
14'd2295:data <=32'hFF5BFFCA;14'd2296:data <=32'hFF5DFFD7;14'd2297:data <=32'hFF5DFFE1;
14'd2298:data <=32'hFF5AFFEC;14'd2299:data <=32'hFF56FFFB;14'd2300:data <=32'hFF52000A;
14'd2301:data <=32'hFF50001D;14'd2302:data <=32'hFF520030;14'd2303:data <=32'hFF550044;
14'd2304:data <=32'hFFC7FFD5;14'd2305:data <=32'hFF9CFFCE;14'd2306:data <=32'hFF78FFE6;
14'd2307:data <=32'hFF770077;14'd2308:data <=32'hFF6300C1;14'd2309:data <=32'hFF8800D6;
14'd2310:data <=32'hFFB300E1;14'd2311:data <=32'hFFDF00E2;14'd2312:data <=32'h000A00D5;
14'd2313:data <=32'h002D00BD;14'd2314:data <=32'h0044009E;14'd2315:data <=32'h004D007C;
14'd2316:data <=32'h004A005F;14'd2317:data <=32'h003E004A;14'd2318:data <=32'h00310040;
14'd2319:data <=32'h0024003F;14'd2320:data <=32'h001D0045;14'd2321:data <=32'h001B004D;
14'd2322:data <=32'h001E0054;14'd2323:data <=32'h0026005B;14'd2324:data <=32'h00300061;
14'd2325:data <=32'h003E0063;14'd2326:data <=32'h004E0063;14'd2327:data <=32'h0063005F;
14'd2328:data <=32'h00770053;14'd2329:data <=32'h00890041;14'd2330:data <=32'h00980027;
14'd2331:data <=32'h009D0007;14'd2332:data <=32'h0097FFE6;14'd2333:data <=32'h0087FFC8;
14'd2334:data <=32'h006CFFB3;14'd2335:data <=32'h004DFFA9;14'd2336:data <=32'h002EFFAB;
14'd2337:data <=32'h0017FFB7;14'd2338:data <=32'h0005FFC9;14'd2339:data <=32'hFFFEFFDF;
14'd2340:data <=32'hFFFEFFF2;14'd2341:data <=32'h00060003;14'd2342:data <=32'h0011000F;
14'd2343:data <=32'h001F0017;14'd2344:data <=32'h002F001B;14'd2345:data <=32'h0040001A;
14'd2346:data <=32'h00520015;14'd2347:data <=32'h0063000B;14'd2348:data <=32'h0073FFFC;
14'd2349:data <=32'h0080FFE8;14'd2350:data <=32'h0086FFCE;14'd2351:data <=32'h0085FFB3;
14'd2352:data <=32'h007FFF99;14'd2353:data <=32'h0072FF82;14'd2354:data <=32'h0063FF6F;
14'd2355:data <=32'h0050FF60;14'd2356:data <=32'h0041FF53;14'd2357:data <=32'h0031FF46;
14'd2358:data <=32'h001FFF37;14'd2359:data <=32'h0009FF27;14'd2360:data <=32'hFFEBFF16;
14'd2361:data <=32'hFFC4FF0A;14'd2362:data <=32'hFF96FF07;14'd2363:data <=32'hFF65FF11;
14'd2364:data <=32'hFF34FF27;14'd2365:data <=32'hFF09FF4C;14'd2366:data <=32'hFEE8FF7A;
14'd2367:data <=32'hFED2FFAF;14'd2368:data <=32'hFFD8FFDE;14'd2369:data <=32'hFFC1FFC3;
14'd2370:data <=32'hFF8EFFAF;14'd2371:data <=32'hFEDEFFF2;14'd2372:data <=32'hFEBB005F;
14'd2373:data <=32'hFEDE009A;14'd2374:data <=32'hFF0F00C8;14'd2375:data <=32'hFF4700E8;
14'd2376:data <=32'hFF8500F5;14'd2377:data <=32'hFFC300F0;14'd2378:data <=32'hFFF500DB;
14'd2379:data <=32'h001A00B9;14'd2380:data <=32'h002E0093;14'd2381:data <=32'h00340070;
14'd2382:data <=32'h002E0053;14'd2383:data <=32'h00230041;14'd2384:data <=32'h00160036;
14'd2385:data <=32'h000B0033;14'd2386:data <=32'h00010033;14'd2387:data <=32'hFFF80037;
14'd2388:data <=32'hFFF4003F;14'd2389:data <=32'hFFF20048;14'd2390:data <=32'hFFF40053;
14'd2391:data <=32'hFFFB0060;14'd2392:data <=32'h0009006A;14'd2393:data <=32'h001C0070;
14'd2394:data <=32'h0031006F;14'd2395:data <=32'h00440065;14'd2396:data <=32'h00540056;
14'd2397:data <=32'h005C0042;14'd2398:data <=32'h005E0030;14'd2399:data <=32'h00590021;
14'd2400:data <=32'h00520017;14'd2401:data <=32'h004A0012;14'd2402:data <=32'h00440011;
14'd2403:data <=32'h00440011;14'd2404:data <=32'h00450010;14'd2405:data <=32'h0048000C;
14'd2406:data <=32'h00490005;14'd2407:data <=32'h0047FFFE;14'd2408:data <=32'h0042FFF9;
14'd2409:data <=32'h003AFFF6;14'd2410:data <=32'h0034FFF8;14'd2411:data <=32'h002FFFFC;
14'd2412:data <=32'h002E0003;14'd2413:data <=32'h0030000A;14'd2414:data <=32'h00370010;
14'd2415:data <=32'h00400015;14'd2416:data <=32'h004C0018;14'd2417:data <=32'h005B0018;
14'd2418:data <=32'h006C0015;14'd2419:data <=32'h00800010;14'd2420:data <=32'h00970002;
14'd2421:data <=32'h00B0FFEC;14'd2422:data <=32'h00C6FFCA;14'd2423:data <=32'h00D3FF9D;
14'd2424:data <=32'h00D5FF67;14'd2425:data <=32'h00C4FF2E;14'd2426:data <=32'h00A2FEF6;
14'd2427:data <=32'h006DFEC9;14'd2428:data <=32'h002CFEAA;14'd2429:data <=32'hFFE5FE9E;
14'd2430:data <=32'hFF9CFEA5;14'd2431:data <=32'hFF59FEBD;14'd2432:data <=32'hFFC0FF67;
14'd2433:data <=32'hFFA5FF53;14'd2434:data <=32'hFF8AFF35;14'd2435:data <=32'hFF46FEEF;
14'd2436:data <=32'hFEECFF4F;14'd2437:data <=32'hFEDAFF89;14'd2438:data <=32'hFED5FFC3;
14'd2439:data <=32'hFEDEFFFD;14'd2440:data <=32'hFEF5002E;14'd2441:data <=32'hFF170054;
14'd2442:data <=32'hFF3A006A;14'd2443:data <=32'hFF5C0075;14'd2444:data <=32'hFF780079;
14'd2445:data <=32'hFF8E0078;14'd2446:data <=32'hFF9D0078;14'd2447:data <=32'hFFAA007A;
14'd2448:data <=32'hFFB8007C;14'd2449:data <=32'hFFC80080;14'd2450:data <=32'hFFD9007F;
14'd2451:data <=32'hFFEB007B;14'd2452:data <=32'hFFFB0072;14'd2453:data <=32'h00060068;
14'd2454:data <=32'h000E005C;14'd2455:data <=32'h00130052;14'd2456:data <=32'h00150049;
14'd2457:data <=32'h00160041;14'd2458:data <=32'h0017003A;14'd2459:data <=32'h00180032;
14'd2460:data <=32'h00130029;14'd2461:data <=32'h000C0022;14'd2462:data <=32'h0003001F;
14'd2463:data <=32'hFFF60022;14'd2464:data <=32'hFFEC002C;14'd2465:data <=32'hFFE6003B;
14'd2466:data <=32'hFFE9004E;14'd2467:data <=32'hFFF30060;14'd2468:data <=32'h0006006D;
14'd2469:data <=32'h001E0072;14'd2470:data <=32'h0036006F;14'd2471:data <=32'h004B0063;
14'd2472:data <=32'h00590052;14'd2473:data <=32'h0060003E;14'd2474:data <=32'h0061002C;
14'd2475:data <=32'h005D001D;14'd2476:data <=32'h00540012;14'd2477:data <=32'h004B000D;
14'd2478:data <=32'h0043000B;14'd2479:data <=32'h003C000D;14'd2480:data <=32'h00370013;
14'd2481:data <=32'h0035001C;14'd2482:data <=32'h00380027;14'd2483:data <=32'h00410035;
14'd2484:data <=32'h00540040;14'd2485:data <=32'h006F0046;14'd2486:data <=32'h00900042;
14'd2487:data <=32'h00B40031;14'd2488:data <=32'h00D30011;14'd2489:data <=32'h00E9FFE4;
14'd2490:data <=32'h00F2FFB0;14'd2491:data <=32'h00EAFF7A;14'd2492:data <=32'h00D2FF47;
14'd2493:data <=32'h00AFFF1E;14'd2494:data <=32'h0083FEFE;14'd2495:data <=32'h0055FEEA;
14'd2496:data <=32'h008DFF0E;14'd2497:data <=32'h0066FED8;14'd2498:data <=32'h0043FEBC;
14'd2499:data <=32'h0044FEFE;14'd2500:data <=32'hFFEFFF28;14'd2501:data <=32'hFFD3FF2E;
14'd2502:data <=32'hFFBCFF39;14'd2503:data <=32'hFFA5FF46;14'd2504:data <=32'hFF95FF55;
14'd2505:data <=32'hFF86FF63;14'd2506:data <=32'hFF79FF6E;14'd2507:data <=32'hFF6BFF79;
14'd2508:data <=32'hFF58FF85;14'd2509:data <=32'hFF43FF95;14'd2510:data <=32'hFF2CFFAF;
14'd2511:data <=32'hFF19FFD1;14'd2512:data <=32'hFF10FFFB;14'd2513:data <=32'hFF130029;
14'd2514:data <=32'hFF240055;14'd2515:data <=32'hFF3F007B;14'd2516:data <=32'hFF640096;
14'd2517:data <=32'hFF8C00A5;14'd2518:data <=32'hFFB400AB;14'd2519:data <=32'hFFD900A7;
14'd2520:data <=32'hFFFA009A;14'd2521:data <=32'h00160088;14'd2522:data <=32'h002C0070;
14'd2523:data <=32'h003A0053;14'd2524:data <=32'h00400033;14'd2525:data <=32'h003B0013;
14'd2526:data <=32'h002AFFF8;14'd2527:data <=32'h0011FFE5;14'd2528:data <=32'hFFF3FFDD;
14'd2529:data <=32'hFFD4FFE2;14'd2530:data <=32'hFFBAFFF3;14'd2531:data <=32'hFFA8000C;
14'd2532:data <=32'hFFA20029;14'd2533:data <=32'hFFA50044;14'd2534:data <=32'hFFB3005C;
14'd2535:data <=32'hFFC4006C;14'd2536:data <=32'hFFD60076;14'd2537:data <=32'hFFE8007C;
14'd2538:data <=32'hFFF7007E;14'd2539:data <=32'h0005007F;14'd2540:data <=32'h0013007F;
14'd2541:data <=32'h001F007F;14'd2542:data <=32'h002E007E;14'd2543:data <=32'h003C007B;
14'd2544:data <=32'h00490075;14'd2545:data <=32'h0055006F;14'd2546:data <=32'h00600068;
14'd2547:data <=32'h006B0063;14'd2548:data <=32'h0076005D;14'd2549:data <=32'h00840058;
14'd2550:data <=32'h0097004E;14'd2551:data <=32'h00AA003F;14'd2552:data <=32'h00BC0029;
14'd2553:data <=32'h00C9000A;14'd2554:data <=32'h00CEFFE8;14'd2555:data <=32'h00C7FFC4;
14'd2556:data <=32'h00B8FFA5;14'd2557:data <=32'h00A1FF8D;14'd2558:data <=32'h0087FF7E;
14'd2559:data <=32'h0070FF79;14'd2560:data <=32'h0124FFCE;14'd2561:data <=32'h0131FF82;
14'd2562:data <=32'h0114FF45;14'd2563:data <=32'h0071FF84;14'd2564:data <=32'h003AFFAE;
14'd2565:data <=32'h003FFFAF;14'd2566:data <=32'h0045FFAB;14'd2567:data <=32'h004BFFA1;
14'd2568:data <=32'h004FFF93;14'd2569:data <=32'h0052FF80;14'd2570:data <=32'h004EFF66;
14'd2571:data <=32'h0040FF4A;14'd2572:data <=32'h0027FF2C;14'd2573:data <=32'h0001FF15;
14'd2574:data <=32'hFFD0FF0A;14'd2575:data <=32'hFF9AFF0D;14'd2576:data <=32'hFF66FF23;
14'd2577:data <=32'hFF39FF48;14'd2578:data <=32'hFF1AFF77;14'd2579:data <=32'hFF0BFFAC;
14'd2580:data <=32'hFF0AFFE1;14'd2581:data <=32'hFF16000F;14'd2582:data <=32'hFF2A0038;
14'd2583:data <=32'hFF470059;14'd2584:data <=32'hFF660072;14'd2585:data <=32'hFF8A0082;
14'd2586:data <=32'hFFB00089;14'd2587:data <=32'hFFD50086;14'd2588:data <=32'hFFF80078;
14'd2589:data <=32'h00120063;14'd2590:data <=32'h00230046;14'd2591:data <=32'h002A0028;
14'd2592:data <=32'h0024000B;14'd2593:data <=32'h0017FFF3;14'd2594:data <=32'h0004FFE5;
14'd2595:data <=32'hFFF0FFDE;14'd2596:data <=32'hFFDDFFDD;14'd2597:data <=32'hFFCDFFE2;
14'd2598:data <=32'hFFBEFFE6;14'd2599:data <=32'hFFB2FFEE;14'd2600:data <=32'hFFA5FFF6;
14'd2601:data <=32'hFF970000;14'd2602:data <=32'hFF88000F;14'd2603:data <=32'hFF7A0024;
14'd2604:data <=32'hFF71003F;14'd2605:data <=32'hFF6F0060;14'd2606:data <=32'hFF760083;
14'd2607:data <=32'hFF8700A7;14'd2608:data <=32'hFFA000C5;14'd2609:data <=32'hFFC100DE;
14'd2610:data <=32'hFFE800EE;14'd2611:data <=32'h001000F8;14'd2612:data <=32'h003C00FA;
14'd2613:data <=32'h006800F3;14'd2614:data <=32'h009500E3;14'd2615:data <=32'h00C000C8;
14'd2616:data <=32'h00E500A2;14'd2617:data <=32'h01000072;14'd2618:data <=32'h010D003C;
14'd2619:data <=32'h010B0003;14'd2620:data <=32'h00F7FFD1;14'd2621:data <=32'h00D7FFA8;
14'd2622:data <=32'h00B0FF90;14'd2623:data <=32'h0088FF86;14'd2624:data <=32'h00B8005E;
14'd2625:data <=32'h00E40040;14'd2626:data <=32'h00FD0004;14'd2627:data <=32'h0093FF90;
14'd2628:data <=32'h004DFFBC;14'd2629:data <=32'h0049FFC6;14'd2630:data <=32'h004BFFCE;
14'd2631:data <=32'h0050FFD2;14'd2632:data <=32'h0059FFD1;14'd2633:data <=32'h0064FFCB;
14'd2634:data <=32'h0070FFBE;14'd2635:data <=32'h007AFFA9;14'd2636:data <=32'h007AFF8B;
14'd2637:data <=32'h006FFF6C;14'd2638:data <=32'h0058FF4E;14'd2639:data <=32'h0035FF3A;
14'd2640:data <=32'h000EFF30;14'd2641:data <=32'hFFE6FF31;14'd2642:data <=32'hFFC3FF40;
14'd2643:data <=32'hFFA6FF55;14'd2644:data <=32'hFF92FF6E;14'd2645:data <=32'hFF85FF86;
14'd2646:data <=32'hFF7EFF9F;14'd2647:data <=32'hFF79FFB5;14'd2648:data <=32'hFF77FFCA;
14'd2649:data <=32'hFF79FFDF;14'd2650:data <=32'hFF7EFFF5;14'd2651:data <=32'hFF870008;
14'd2652:data <=32'hFF950017;14'd2653:data <=32'hFFA50022;14'd2654:data <=32'hFFB60028;
14'd2655:data <=32'hFFC50028;14'd2656:data <=32'hFFD20026;14'd2657:data <=32'hFFDC0021;
14'd2658:data <=32'hFFE4001D;14'd2659:data <=32'hFFEC0019;14'd2660:data <=32'hFFF30012;
14'd2661:data <=32'hFFFB0009;14'd2662:data <=32'h0003FFFC;14'd2663:data <=32'h0006FFE9;
14'd2664:data <=32'h0000FFD3;14'd2665:data <=32'hFFF2FFBB;14'd2666:data <=32'hFFD8FFA9;
14'd2667:data <=32'hFFB5FF9E;14'd2668:data <=32'hFF8FFFA1;14'd2669:data <=32'hFF66FFB2;
14'd2670:data <=32'hFF43FFCF;14'd2671:data <=32'hFF28FFF7;14'd2672:data <=32'hFF180027;
14'd2673:data <=32'hFF150059;14'd2674:data <=32'hFF20008E;14'd2675:data <=32'hFF3400BE;
14'd2676:data <=32'hFF5500EB;14'd2677:data <=32'hFF800110;14'd2678:data <=32'hFFB5012C;
14'd2679:data <=32'hFFF2013B;14'd2680:data <=32'h0031013B;14'd2681:data <=32'h006E0129;
14'd2682:data <=32'h00A50106;14'd2683:data <=32'h00CE00D9;14'd2684:data <=32'h00E800A4;
14'd2685:data <=32'h00F0006E;14'd2686:data <=32'h00E9003F;14'd2687:data <=32'h00D9001B;
14'd2688:data <=32'h008B004A;14'd2689:data <=32'h009D0044;14'd2690:data <=32'h00BE0039;
14'd2691:data <=32'h00FB0025;14'd2692:data <=32'h00C30030;14'd2693:data <=32'h00C6001A;
14'd2694:data <=32'h00C70002;14'd2695:data <=32'h00C4FFE9;14'd2696:data <=32'h00BDFFD2;
14'd2697:data <=32'h00B3FFBD;14'd2698:data <=32'h00A9FFAA;14'd2699:data <=32'h009EFF96;
14'd2700:data <=32'h008EFF82;14'd2701:data <=32'h007AFF6E;14'd2702:data <=32'h005FFF5F;
14'd2703:data <=32'h003FFF57;14'd2704:data <=32'h001DFF58;14'd2705:data <=32'hFFFFFF64;
14'd2706:data <=32'hFFE7FF77;14'd2707:data <=32'hFFDAFF8F;14'd2708:data <=32'hFFD7FFA8;
14'd2709:data <=32'hFFDBFFBA;14'd2710:data <=32'hFFE6FFC4;14'd2711:data <=32'hFFF0FFC8;
14'd2712:data <=32'hFFF6FFC5;14'd2713:data <=32'hFFF9FFBF;14'd2714:data <=32'hFFF7FFBA;
14'd2715:data <=32'hFFF2FFB5;14'd2716:data <=32'hFFEBFFB3;14'd2717:data <=32'hFFE3FFB1;
14'd2718:data <=32'hFFDAFFB2;14'd2719:data <=32'hFFD1FFB4;14'd2720:data <=32'hFFC6FFB9;
14'd2721:data <=32'hFFBDFFC2;14'd2722:data <=32'hFFB4FFCE;14'd2723:data <=32'hFFB0FFDF;
14'd2724:data <=32'hFFB3FFF0;14'd2725:data <=32'hFFBEFFFE;14'd2726:data <=32'hFFCF0008;
14'd2727:data <=32'hFFE40008;14'd2728:data <=32'hFFF5FFFF;14'd2729:data <=32'h0003FFEB;
14'd2730:data <=32'h0005FFD4;14'd2731:data <=32'hFFFDFFB9;14'd2732:data <=32'hFFEAFFA4;
14'd2733:data <=32'hFFCFFF95;14'd2734:data <=32'hFFAEFF92;14'd2735:data <=32'hFF8EFF97;
14'd2736:data <=32'hFF6FFFA6;14'd2737:data <=32'hFF55FFBC;14'd2738:data <=32'hFF3FFFD8;
14'd2739:data <=32'hFF30FFF8;14'd2740:data <=32'hFF27001C;14'd2741:data <=32'hFF240043;
14'd2742:data <=32'hFF2A006A;14'd2743:data <=32'hFF3A0092;14'd2744:data <=32'hFF5400B5;
14'd2745:data <=32'hFF7500D1;14'd2746:data <=32'hFF9B00E2;14'd2747:data <=32'hFFBF00E9;
14'd2748:data <=32'hFFE100E9;14'd2749:data <=32'hFFFE00E4;14'd2750:data <=32'h001500DE;
14'd2751:data <=32'h002900DB;14'd2752:data <=32'h008700AC;14'd2753:data <=32'h0099009D;
14'd2754:data <=32'h009E009C;14'd2755:data <=32'h005E0103;14'd2756:data <=32'h00550122;
14'd2757:data <=32'h008C0116;14'd2758:data <=32'h00C000FB;14'd2759:data <=32'h00EE00D3;
14'd2760:data <=32'h010E00A4;14'd2761:data <=32'h0124006E;14'd2762:data <=32'h01300037;
14'd2763:data <=32'h012FFFFE;14'd2764:data <=32'h0122FFC7;14'd2765:data <=32'h0108FF92;
14'd2766:data <=32'h00E3FF65;14'd2767:data <=32'h00B2FF43;14'd2768:data <=32'h007BFF32;
14'd2769:data <=32'h0043FF33;14'd2770:data <=32'h0010FF43;14'd2771:data <=32'hFFE9FF61;
14'd2772:data <=32'hFFD3FF87;14'd2773:data <=32'hFFCAFFAD;14'd2774:data <=32'hFFCFFFCC;
14'd2775:data <=32'hFFDCFFE5;14'd2776:data <=32'hFFEEFFF4;14'd2777:data <=32'h0000FFFA;
14'd2778:data <=32'h0011FFFA;14'd2779:data <=32'h001EFFF7;14'd2780:data <=32'h002AFFEF;
14'd2781:data <=32'h0032FFE4;14'd2782:data <=32'h0037FFD6;14'd2783:data <=32'h0038FFC7;
14'd2784:data <=32'h0034FFB7;14'd2785:data <=32'h002AFFAA;14'd2786:data <=32'h001BFFA0;
14'd2787:data <=32'h000BFF9C;14'd2788:data <=32'hFFFCFF9E;14'd2789:data <=32'hFFF1FFA4;
14'd2790:data <=32'hFFEBFFAC;14'd2791:data <=32'hFFE8FFB2;14'd2792:data <=32'hFFEAFFB4;
14'd2793:data <=32'hFFEBFFB2;14'd2794:data <=32'hFFE9FFAB;14'd2795:data <=32'hFFE3FFA3;
14'd2796:data <=32'hFFD6FF9D;14'd2797:data <=32'hFFC6FF9D;14'd2798:data <=32'hFFB4FFA0;
14'd2799:data <=32'hFFA5FFA9;14'd2800:data <=32'hFF99FFB6;14'd2801:data <=32'hFF92FFC3;
14'd2802:data <=32'hFF8FFFCF;14'd2803:data <=32'hFF8DFFD9;14'd2804:data <=32'hFF8DFFE0;
14'd2805:data <=32'hFF8AFFE7;14'd2806:data <=32'hFF87FFED;14'd2807:data <=32'hFF82FFF4;
14'd2808:data <=32'hFF7CFFFD;14'd2809:data <=32'hFF780006;14'd2810:data <=32'hFF73000E;
14'd2811:data <=32'hFF6C0017;14'd2812:data <=32'hFF630022;14'd2813:data <=32'hFF560031;
14'd2814:data <=32'hFF480049;14'd2815:data <=32'hFF3D006A;14'd2816:data <=32'hFFBA00D5;
14'd2817:data <=32'hFFD000E7;14'd2818:data <=32'hFFD900E0;14'd2819:data <=32'hFF5D00B7;
14'd2820:data <=32'hFF430107;14'd2821:data <=32'hFF790132;14'd2822:data <=32'hFFB7014E;
14'd2823:data <=32'hFFFA0156;14'd2824:data <=32'h003D0150;14'd2825:data <=32'h007A013C;
14'd2826:data <=32'h00B2011D;14'd2827:data <=32'h00E100F1;14'd2828:data <=32'h010500BC;
14'd2829:data <=32'h011D0081;14'd2830:data <=32'h01240041;14'd2831:data <=32'h011B0003;
14'd2832:data <=32'h0101FFCC;14'd2833:data <=32'h00DBFFA2;14'd2834:data <=32'h00AEFF88;
14'd2835:data <=32'h0081FF7D;14'd2836:data <=32'h0059FF80;14'd2837:data <=32'h003AFF8B;
14'd2838:data <=32'h0024FF9A;14'd2839:data <=32'h0016FFA9;14'd2840:data <=32'h000BFFB7;
14'd2841:data <=32'h0005FFC4;14'd2842:data <=32'hFFFFFFD0;14'd2843:data <=32'hFFFDFFDD;
14'd2844:data <=32'hFFFDFFEC;14'd2845:data <=32'h0000FFF9;14'd2846:data <=32'h000B0004;
14'd2847:data <=32'h0017000C;14'd2848:data <=32'h0027000E;14'd2849:data <=32'h0035000B;
14'd2850:data <=32'h00420004;14'd2851:data <=32'h004DFFFB;14'd2852:data <=32'h0055FFEF;
14'd2853:data <=32'h005BFFE2;14'd2854:data <=32'h0063FFD4;14'd2855:data <=32'h0067FFC2;
14'd2856:data <=32'h0068FFAC;14'd2857:data <=32'h0065FF94;14'd2858:data <=32'h0059FF79;
14'd2859:data <=32'h0044FF5F;14'd2860:data <=32'h0026FF4B;14'd2861:data <=32'h0002FF41;
14'd2862:data <=32'hFFDBFF42;14'd2863:data <=32'hFFB7FF4E;14'd2864:data <=32'hFF9AFF65;
14'd2865:data <=32'hFF86FF81;14'd2866:data <=32'hFF7DFF9F;14'd2867:data <=32'hFF7EFFBC;
14'd2868:data <=32'hFF85FFD0;14'd2869:data <=32'hFF8FFFE1;14'd2870:data <=32'hFF9BFFE9;
14'd2871:data <=32'hFFA8FFEE;14'd2872:data <=32'hFFB1FFEC;14'd2873:data <=32'hFFB9FFE6;
14'd2874:data <=32'hFFBCFFDB;14'd2875:data <=32'hFFB9FFCF;14'd2876:data <=32'hFFADFFC0;
14'd2877:data <=32'hFF97FFB5;14'd2878:data <=32'hFF77FFB1;14'd2879:data <=32'hFF53FFBB;
14'd2880:data <=32'hFF51FFF9;14'd2881:data <=32'hFF310012;14'd2882:data <=32'hFF2F002A;
14'd2883:data <=32'hFF50000D;14'd2884:data <=32'hFF130055;14'd2885:data <=32'hFF220081;
14'd2886:data <=32'hFF3C00A8;14'd2887:data <=32'hFF5E00C6;14'd2888:data <=32'hFF8200DA;
14'd2889:data <=32'hFFA700E8;14'd2890:data <=32'hFFCC00EF;14'd2891:data <=32'hFFF200F0;
14'd2892:data <=32'h001800EB;14'd2893:data <=32'h003B00DE;14'd2894:data <=32'h005B00C9;
14'd2895:data <=32'h007300AF;14'd2896:data <=32'h00830091;14'd2897:data <=32'h008B0075;
14'd2898:data <=32'h008C005D;14'd2899:data <=32'h008A004A;14'd2900:data <=32'h0087003A;
14'd2901:data <=32'h0087002D;14'd2902:data <=32'h00890020;14'd2903:data <=32'h008B000E;
14'd2904:data <=32'h008AFFF9;14'd2905:data <=32'h0083FFE2;14'd2906:data <=32'h0073FFCD;
14'd2907:data <=32'h005EFFBD;14'd2908:data <=32'h0044FFB5;14'd2909:data <=32'h0029FFB6;
14'd2910:data <=32'h0011FFBF;14'd2911:data <=32'h0000FFD1;14'd2912:data <=32'hFFF5FFE5;
14'd2913:data <=32'hFFF2FFFA;14'd2914:data <=32'hFFF5000F;14'd2915:data <=32'hFFFE0023;
14'd2916:data <=32'h000D0034;14'd2917:data <=32'h00230041;14'd2918:data <=32'h003D0047;
14'd2919:data <=32'h005B0046;14'd2920:data <=32'h007B003A;14'd2921:data <=32'h009A0023;
14'd2922:data <=32'h00B00001;14'd2923:data <=32'h00BBFFD8;14'd2924:data <=32'h00B8FFAB;
14'd2925:data <=32'h00A9FF81;14'd2926:data <=32'h008DFF5E;14'd2927:data <=32'h0069FF46;
14'd2928:data <=32'h0042FF3A;14'd2929:data <=32'h001FFF3A;14'd2930:data <=32'h0000FF40;
14'd2931:data <=32'hFFE7FF4C;14'd2932:data <=32'hFFD5FF58;14'd2933:data <=32'hFFC6FF66;
14'd2934:data <=32'hFFBAFF71;14'd2935:data <=32'hFFB1FF7C;14'd2936:data <=32'hFFA9FF87;
14'd2937:data <=32'hFFA3FF91;14'd2938:data <=32'hFFA0FF99;14'd2939:data <=32'hFF9CFF9D;
14'd2940:data <=32'hFF97FF9F;14'd2941:data <=32'hFF8EFF9F;14'd2942:data <=32'hFF7EFF9F;
14'd2943:data <=32'hFF69FFA4;14'd2944:data <=32'hFFEAFF7B;14'd2945:data <=32'hFFB5FF5F;
14'd2946:data <=32'hFF81FF6A;14'd2947:data <=32'hFF55FFF1;14'd2948:data <=32'hFF1E002F;
14'd2949:data <=32'hFF340053;14'd2950:data <=32'hFF51006D;14'd2951:data <=32'hFF73007B;
14'd2952:data <=32'hFF90007F;14'd2953:data <=32'hFFA9007B;14'd2954:data <=32'hFFBA0075;
14'd2955:data <=32'hFFC5006D;14'd2956:data <=32'hFFCD0068;14'd2957:data <=32'hFFD30063;
14'd2958:data <=32'hFFD60060;14'd2959:data <=32'hFFD7005E;14'd2960:data <=32'hFFD7005E;
14'd2961:data <=32'hFFD50061;14'd2962:data <=32'hFFD4006B;14'd2963:data <=32'hFFD70078;
14'd2964:data <=32'hFFE10089;14'd2965:data <=32'hFFF3009A;14'd2966:data <=32'h000F00A6;
14'd2967:data <=32'h003000A8;14'd2968:data <=32'h0054009D;14'd2969:data <=32'h00720086;
14'd2970:data <=32'h00880069;14'd2971:data <=32'h00920045;14'd2972:data <=32'h00900021;
14'd2973:data <=32'h00840003;14'd2974:data <=32'h0071FFEC;14'd2975:data <=32'h0059FFDD;
14'd2976:data <=32'h0043FFD6;14'd2977:data <=32'h002CFFD5;14'd2978:data <=32'h0017FFDC;
14'd2979:data <=32'h0006FFE7;14'd2980:data <=32'hFFF8FFF8;14'd2981:data <=32'hFFF1000D;
14'd2982:data <=32'hFFF10025;14'd2983:data <=32'hFFFB003D;14'd2984:data <=32'h000D0050;
14'd2985:data <=32'h0027005E;14'd2986:data <=32'h00450061;14'd2987:data <=32'h0062005A;
14'd2988:data <=32'h007D004A;14'd2989:data <=32'h00900035;14'd2990:data <=32'h009D001C;
14'd2991:data <=32'h00A30005;14'd2992:data <=32'h00A4FFEF;14'd2993:data <=32'h00A5FFDB;
14'd2994:data <=32'h00A6FFC8;14'd2995:data <=32'h00A7FFB3;14'd2996:data <=32'h00A8FF9C;
14'd2997:data <=32'h00A4FF7E;14'd2998:data <=32'h0099FF60;14'd2999:data <=32'h0086FF40;
14'd3000:data <=32'h006BFF24;14'd3001:data <=32'h004AFF0D;14'd3002:data <=32'h0024FEFE;
14'd3003:data <=32'hFFFCFEF6;14'd3004:data <=32'hFFD2FEF5;14'd3005:data <=32'hFFA7FEF9;
14'd3006:data <=32'hFF7CFF06;14'd3007:data <=32'hFF4FFF1B;14'd3008:data <=32'h002BFFAE;
14'd3009:data <=32'h001AFF7B;14'd3010:data <=32'hFFE8FF50;14'd3011:data <=32'hFF20FF5D;
14'd3012:data <=32'hFED4FFB3;14'd3013:data <=32'hFEDFFFF4;14'd3014:data <=32'hFEFA0029;
14'd3015:data <=32'hFF210054;14'd3016:data <=32'hFF4C006B;14'd3017:data <=32'hFF770074;
14'd3018:data <=32'hFF9A0071;14'd3019:data <=32'hFFB60067;14'd3020:data <=32'hFFCA005A;
14'd3021:data <=32'hFFD9004A;14'd3022:data <=32'hFFDF003A;14'd3023:data <=32'hFFDF002A;
14'd3024:data <=32'hFFD9001D;14'd3025:data <=32'hFFCD0014;14'd3026:data <=32'hFFBC0012;
14'd3027:data <=32'hFFAB001B;14'd3028:data <=32'hFF9E002C;14'd3029:data <=32'hFF980044;
14'd3030:data <=32'hFF9D005F;14'd3031:data <=32'hFFAD0077;14'd3032:data <=32'hFFC50089;
14'd3033:data <=32'hFFE20092;14'd3034:data <=32'hFFFD008F;14'd3035:data <=32'h00150085;
14'd3036:data <=32'h00260076;14'd3037:data <=32'h00310067;14'd3038:data <=32'h00380059;
14'd3039:data <=32'h003A004D;14'd3040:data <=32'h003B0041;14'd3041:data <=32'h003D0037;
14'd3042:data <=32'h003C002D;14'd3043:data <=32'h00380023;14'd3044:data <=32'h0033001B;
14'd3045:data <=32'h002B0015;14'd3046:data <=32'h00210013;14'd3047:data <=32'h00190016;
14'd3048:data <=32'h0013001B;14'd3049:data <=32'h00100023;14'd3050:data <=32'h0010002B;
14'd3051:data <=32'h00120031;14'd3052:data <=32'h00140037;14'd3053:data <=32'h0018003D;
14'd3054:data <=32'h001C0045;14'd3055:data <=32'h0021004F;14'd3056:data <=32'h002A005D;
14'd3057:data <=32'h003A006C;14'd3058:data <=32'h00540079;14'd3059:data <=32'h0077007F;
14'd3060:data <=32'h00A1007B;14'd3061:data <=32'h00CC0067;14'd3062:data <=32'h00F40043;
14'd3063:data <=32'h01130015;14'd3064:data <=32'h0124FFDD;14'd3065:data <=32'h0128FFA0;
14'd3066:data <=32'h011BFF62;14'd3067:data <=32'h0100FF29;14'd3068:data <=32'h00DBFEF5;
14'd3069:data <=32'h00A8FEC9;14'd3070:data <=32'h006CFEA8;14'd3071:data <=32'h0028FE94;
14'd3072:data <=32'h003EFF70;14'd3073:data <=32'h0032FF48;14'd3074:data <=32'h0023FF16;
14'd3075:data <=32'hFFE7FEAE;14'd3076:data <=32'hFF6CFEE4;14'd3077:data <=32'hFF46FF14;
14'd3078:data <=32'hFF30FF49;14'd3079:data <=32'hFF29FF7B;14'd3080:data <=32'hFF2EFFA3;
14'd3081:data <=32'hFF39FFC5;14'd3082:data <=32'hFF45FFDE;14'd3083:data <=32'hFF51FFF2;
14'd3084:data <=32'hFF5D0004;14'd3085:data <=32'hFF6A0013;14'd3086:data <=32'hFF780020;
14'd3087:data <=32'hFF860028;14'd3088:data <=32'hFF94002D;14'd3089:data <=32'hFF9F002E;
14'd3090:data <=32'hFFA6002D;14'd3091:data <=32'hFFAA002D;14'd3092:data <=32'hFFAC0031;
14'd3093:data <=32'hFFAF0037;14'd3094:data <=32'hFFB5003F;14'd3095:data <=32'hFFBF0047;
14'd3096:data <=32'hFFCD004A;14'd3097:data <=32'hFFDB0048;14'd3098:data <=32'hFFE60041;
14'd3099:data <=32'hFFEB0036;14'd3100:data <=32'hFFEB002B;14'd3101:data <=32'hFFE40024;
14'd3102:data <=32'hFFDB0023;14'd3103:data <=32'hFFD10027;14'd3104:data <=32'hFFCA0031;
14'd3105:data <=32'hFFCA003F;14'd3106:data <=32'hFFCF004D;14'd3107:data <=32'hFFD90057;
14'd3108:data <=32'hFFE6005E;14'd3109:data <=32'hFFF20061;14'd3110:data <=32'h00000061;
14'd3111:data <=32'h000C005E;14'd3112:data <=32'h00170058;14'd3113:data <=32'h001E0051;
14'd3114:data <=32'h00250047;14'd3115:data <=32'h0028003D;14'd3116:data <=32'h00260032;
14'd3117:data <=32'h001E0028;14'd3118:data <=32'h00120023;14'd3119:data <=32'h00020025;
14'd3120:data <=32'hFFF30032;14'd3121:data <=32'hFFE90048;14'd3122:data <=32'hFFEA0065;
14'd3123:data <=32'hFFF80085;14'd3124:data <=32'h001300A0;14'd3125:data <=32'h003B00B4;
14'd3126:data <=32'h006900BB;14'd3127:data <=32'h009B00B1;14'd3128:data <=32'h00C7009A;
14'd3129:data <=32'h00EE0078;14'd3130:data <=32'h010C004C;14'd3131:data <=32'h0120001C;
14'd3132:data <=32'h0129FFE7;14'd3133:data <=32'h0128FFAF;14'd3134:data <=32'h011AFF78;
14'd3135:data <=32'h0101FF43;14'd3136:data <=32'h00FDFF7D;14'd3137:data <=32'h00F6FF39;
14'd3138:data <=32'h00E6FF0E;14'd3139:data <=32'h00D9FF36;14'd3140:data <=32'h0075FF38;
14'd3141:data <=32'h0058FF34;14'd3142:data <=32'h0041FF33;14'd3143:data <=32'h002CFF34;
14'd3144:data <=32'h001BFF31;14'd3145:data <=32'h0008FF2B;14'd3146:data <=32'hFFEFFF25;
14'd3147:data <=32'hFFD1FF22;14'd3148:data <=32'hFFAFFF26;14'd3149:data <=32'hFF8BFF35;
14'd3150:data <=32'hFF6AFF4B;14'd3151:data <=32'hFF51FF69;14'd3152:data <=32'hFF3DFF8B;
14'd3153:data <=32'hFF34FFAF;14'd3154:data <=32'hFF30FFD5;14'd3155:data <=32'hFF34FFF7;
14'd3156:data <=32'hFF3E0019;14'd3157:data <=32'hFF50003A;14'd3158:data <=32'hFF690055;
14'd3159:data <=32'hFF88006A;14'd3160:data <=32'hFFAE0074;14'd3161:data <=32'hFFD40073;
14'd3162:data <=32'hFFF70064;14'd3163:data <=32'h0010004A;14'd3164:data <=32'h001C002B;
14'd3165:data <=32'h001D000B;14'd3166:data <=32'h000FFFF0;14'd3167:data <=32'hFFFBFFDE;
14'd3168:data <=32'hFFE2FFD6;14'd3169:data <=32'hFFCAFFD8;14'd3170:data <=32'hFFB6FFE1;
14'd3171:data <=32'hFFA7FFF0;14'd3172:data <=32'hFF9D0000;14'd3173:data <=32'hFF980013;
14'd3174:data <=32'hFF970025;14'd3175:data <=32'hFF990037;14'd3176:data <=32'hFFA00048;
14'd3177:data <=32'hFFAA0057;14'd3178:data <=32'hFFB70062;14'd3179:data <=32'hFFC6006A;
14'd3180:data <=32'hFFD5006D;14'd3181:data <=32'hFFE2006B;14'd3182:data <=32'hFFEA0067;
14'd3183:data <=32'hFFED0064;14'd3184:data <=32'hFFEC0064;14'd3185:data <=32'hFFEB006A;
14'd3186:data <=32'hFFEC0076;14'd3187:data <=32'hFFF20086;14'd3188:data <=32'h00020097;
14'd3189:data <=32'h001900A3;14'd3190:data <=32'h003600A9;14'd3191:data <=32'h005500A6;
14'd3192:data <=32'h0072009A;14'd3193:data <=32'h008A0088;14'd3194:data <=32'h009C0072;
14'd3195:data <=32'h00A9005C;14'd3196:data <=32'h00B10047;14'd3197:data <=32'h00B70030;
14'd3198:data <=32'h00BC001A;14'd3199:data <=32'h00BD0004;14'd3200:data <=32'h01320074;
14'd3201:data <=32'h01610031;14'd3202:data <=32'h0161FFEE;14'd3203:data <=32'h00BBFFF5;
14'd3204:data <=32'h00780001;14'd3205:data <=32'h00820003;14'd3206:data <=32'h00910000;
14'd3207:data <=32'h00A5FFF5;14'd3208:data <=32'h00BAFFDF;14'd3209:data <=32'h00C9FFBD;
14'd3210:data <=32'h00CFFF91;14'd3211:data <=32'h00C5FF61;14'd3212:data <=32'h00AAFF33;
14'd3213:data <=32'h0082FF0E;14'd3214:data <=32'h0051FEF4;14'd3215:data <=32'h001BFEEA;
14'd3216:data <=32'hFFE6FEEC;14'd3217:data <=32'hFFB3FEFA;14'd3218:data <=32'hFF86FF12;
14'd3219:data <=32'hFF5FFF33;14'd3220:data <=32'hFF42FF5C;14'd3221:data <=32'hFF2DFF8C;
14'd3222:data <=32'hFF26FFBF;14'd3223:data <=32'hFF2DFFF1;14'd3224:data <=32'hFF43001F;
14'd3225:data <=32'hFF640043;14'd3226:data <=32'hFF8C0058;14'd3227:data <=32'hFFB6005E;
14'd3228:data <=32'hFFDB0056;14'd3229:data <=32'hFFF90044;14'd3230:data <=32'h000B002D;
14'd3231:data <=32'h00130015;14'd3232:data <=32'h00140000;14'd3233:data <=32'h000FFFEE;
14'd3234:data <=32'h0007FFDE;14'd3235:data <=32'hFFFEFFD1;14'd3236:data <=32'hFFF2FFC6;
14'd3237:data <=32'hFFE4FFBE;14'd3238:data <=32'hFFD3FFB7;14'd3239:data <=32'hFFBFFFB4;
14'd3240:data <=32'hFFA9FFB6;14'd3241:data <=32'hFF92FFC0;14'd3242:data <=32'hFF7DFFCF;
14'd3243:data <=32'hFF6CFFE3;14'd3244:data <=32'hFF5FFFFA;14'd3245:data <=32'hFF570011;
14'd3246:data <=32'hFF53002C;14'd3247:data <=32'hFF510047;14'd3248:data <=32'hFF530064;
14'd3249:data <=32'hFF5B0084;14'd3250:data <=32'hFF6900A7;14'd3251:data <=32'hFF8200C7;
14'd3252:data <=32'hFFA400E4;14'd3253:data <=32'hFFCF00F9;14'd3254:data <=32'h00000100;
14'd3255:data <=32'h003300FA;14'd3256:data <=32'h006000E5;14'd3257:data <=32'h008400C5;
14'd3258:data <=32'h009C009F;14'd3259:data <=32'h00A60078;14'd3260:data <=32'h00A60056;
14'd3261:data <=32'h009F0039;14'd3262:data <=32'h00920023;14'd3263:data <=32'h00840013;
14'd3264:data <=32'h006F00DD;14'd3265:data <=32'h00AB00D3;14'd3266:data <=32'h00DA00A2;
14'd3267:data <=32'h0095000E;14'd3268:data <=32'h0045001F;14'd3269:data <=32'h00430030;
14'd3270:data <=32'h004D0040;14'd3271:data <=32'h005F004C;14'd3272:data <=32'h007D0051;
14'd3273:data <=32'h009F0046;14'd3274:data <=32'h00BD002D;14'd3275:data <=32'h00D1000A;
14'd3276:data <=32'h00DBFFDF;14'd3277:data <=32'h00D7FFB3;14'd3278:data <=32'h00C6FF8B;
14'd3279:data <=32'h00AEFF6A;14'd3280:data <=32'h008FFF50;14'd3281:data <=32'h006EFF3E;
14'd3282:data <=32'h004BFF32;14'd3283:data <=32'h0027FF2E;14'd3284:data <=32'h0003FF2F;
14'd3285:data <=32'hFFDFFF3A;14'd3286:data <=32'hFFBEFF4C;14'd3287:data <=32'hFFA5FF66;
14'd3288:data <=32'hFF95FF85;14'd3289:data <=32'hFF8EFFA4;14'd3290:data <=32'hFF90FFC1;
14'd3291:data <=32'hFF99FFD7;14'd3292:data <=32'hFFA5FFE8;14'd3293:data <=32'hFFB2FFF3;
14'd3294:data <=32'hFFBCFFF9;14'd3295:data <=32'hFFC4FFFF;14'd3296:data <=32'hFFCC0004;
14'd3297:data <=32'hFFD6000B;14'd3298:data <=32'hFFE3000F;14'd3299:data <=32'hFFF30011;
14'd3300:data <=32'h0006000B;14'd3301:data <=32'h0017FFFE;14'd3302:data <=32'h0025FFE9;
14'd3303:data <=32'h0029FFCF;14'd3304:data <=32'h0024FFB2;14'd3305:data <=32'h0016FF97;
14'd3306:data <=32'hFFFFFF80;14'd3307:data <=32'hFFE1FF70;14'd3308:data <=32'hFFBDFF67;
14'd3309:data <=32'hFF97FF66;14'd3310:data <=32'hFF6FFF70;14'd3311:data <=32'hFF47FF82;
14'd3312:data <=32'hFF22FF9F;14'd3313:data <=32'hFF02FFC7;14'd3314:data <=32'hFEEBFFFA;
14'd3315:data <=32'hFEE20035;14'd3316:data <=32'hFEE80072;14'd3317:data <=32'hFF0100AF;
14'd3318:data <=32'hFF2B00E2;14'd3319:data <=32'hFF600105;14'd3320:data <=32'hFF9C0118;
14'd3321:data <=32'hFFD5011A;14'd3322:data <=32'h0009010C;14'd3323:data <=32'h003400F5;
14'd3324:data <=32'h005200D9;14'd3325:data <=32'h006800BB;14'd3326:data <=32'h0075009F;
14'd3327:data <=32'h007B0084;14'd3328:data <=32'h00230091;14'd3329:data <=32'h00370099;
14'd3330:data <=32'h005E009D;14'd3331:data <=32'h00A3008E;14'd3332:data <=32'h00650086;
14'd3333:data <=32'h006B007E;14'd3334:data <=32'h00750078;14'd3335:data <=32'h00810071;
14'd3336:data <=32'h00900069;14'd3337:data <=32'h00A50059;14'd3338:data <=32'h00B50041;
14'd3339:data <=32'h00C00022;14'd3340:data <=32'h00C10000;14'd3341:data <=32'h00B8FFDF;
14'd3342:data <=32'h00A5FFC5;14'd3343:data <=32'h008FFFB3;14'd3344:data <=32'h0078FFA9;
14'd3345:data <=32'h0064FFA6;14'd3346:data <=32'h0054FFA7;14'd3347:data <=32'h0048FFA9;
14'd3348:data <=32'h003FFFAB;14'd3349:data <=32'h0036FFAC;14'd3350:data <=32'h002EFFAD;
14'd3351:data <=32'h0028FFB0;14'd3352:data <=32'h0022FFB3;14'd3353:data <=32'h0020FFB6;
14'd3354:data <=32'h0021FFB5;14'd3355:data <=32'h0020FFB2;14'd3356:data <=32'h001DFFAB;
14'd3357:data <=32'h0015FFA3;14'd3358:data <=32'h0008FF9C;14'd3359:data <=32'hFFF8FF99;
14'd3360:data <=32'hFFE4FF9E;14'd3361:data <=32'hFFD3FFAB;14'd3362:data <=32'hFFC8FFBF;
14'd3363:data <=32'hFFC6FFD6;14'd3364:data <=32'hFFCDFFEB;14'd3365:data <=32'hFFDFFFFB;
14'd3366:data <=32'hFFF40002;14'd3367:data <=32'h000B0000;14'd3368:data <=32'h001FFFF4;
14'd3369:data <=32'h002EFFE1;14'd3370:data <=32'h0035FFC9;14'd3371:data <=32'h0035FFB0;
14'd3372:data <=32'h002CFF95;14'd3373:data <=32'h001EFF7B;14'd3374:data <=32'h0006FF65;
14'd3375:data <=32'hFFE9FF53;14'd3376:data <=32'hFFC2FF48;14'd3377:data <=32'hFF9AFF47;
14'd3378:data <=32'hFF6CFF52;14'd3379:data <=32'hFF42FF6A;14'd3380:data <=32'hFF20FF8D;
14'd3381:data <=32'hFF08FFBA;14'd3382:data <=32'hFEFEFFEA;14'd3383:data <=32'hFF010018;
14'd3384:data <=32'hFF0F0041;14'd3385:data <=32'hFF220061;14'd3386:data <=32'hFF37007A;
14'd3387:data <=32'hFF4B008D;14'd3388:data <=32'hFF5E009E;14'd3389:data <=32'hFF7000AE;
14'd3390:data <=32'hFF8400C0;14'd3391:data <=32'hFF9C00CF;14'd3392:data <=32'h000C00B4;
14'd3393:data <=32'h001E00AF;14'd3394:data <=32'h001F00B2;14'd3395:data <=32'hFFCB0103;
14'd3396:data <=32'hFFB10119;14'd3397:data <=32'hFFDF0127;14'd3398:data <=32'h0010012D;
14'd3399:data <=32'h00430128;14'd3400:data <=32'h00780118;14'd3401:data <=32'h00AB00FD;
14'd3402:data <=32'h00D700D3;14'd3403:data <=32'h00F7009E;14'd3404:data <=32'h01060060;
14'd3405:data <=32'h01030024;14'd3406:data <=32'h00EFFFEE;14'd3407:data <=32'h00CDFFC4;
14'd3408:data <=32'h00A5FFA9;14'd3409:data <=32'h007CFF9D;14'd3410:data <=32'h0058FF9E;
14'd3411:data <=32'h003BFFA7;14'd3412:data <=32'h0024FFB5;14'd3413:data <=32'h0015FFC7;
14'd3414:data <=32'h000CFFD8;14'd3415:data <=32'h000AFFEB;14'd3416:data <=32'h000EFFFB;
14'd3417:data <=32'h0018000A;14'd3418:data <=32'h00290013;14'd3419:data <=32'h003A0014;
14'd3420:data <=32'h004E000C;14'd3421:data <=32'h005CFFFD;14'd3422:data <=32'h0063FFE8;
14'd3423:data <=32'h0061FFD2;14'd3424:data <=32'h0056FFBF;14'd3425:data <=32'h0046FFB3;
14'd3426:data <=32'h0035FFAE;14'd3427:data <=32'h0025FFB0;14'd3428:data <=32'h001AFFB6;
14'd3429:data <=32'h0017FFBE;14'd3430:data <=32'h0017FFC4;14'd3431:data <=32'h001AFFC6;
14'd3432:data <=32'h001EFFC5;14'd3433:data <=32'h0020FFC0;14'd3434:data <=32'h0021FFBA;
14'd3435:data <=32'h001DFFB3;14'd3436:data <=32'h001AFFAC;14'd3437:data <=32'h0016FFA6;
14'd3438:data <=32'h0011FF9F;14'd3439:data <=32'h000BFF97;14'd3440:data <=32'h0003FF8F;
14'd3441:data <=32'hFFF8FF87;14'd3442:data <=32'hFFE9FF81;14'd3443:data <=32'hFFD8FF7E;
14'd3444:data <=32'hFFC7FF80;14'd3445:data <=32'hFFB7FF86;14'd3446:data <=32'hFFABFF8C;
14'd3447:data <=32'hFFA1FF93;14'd3448:data <=32'hFF9AFF96;14'd3449:data <=32'hFF90FF97;
14'd3450:data <=32'hFF81FF95;14'd3451:data <=32'hFF6AFF94;14'd3452:data <=32'hFF4EFF99;
14'd3453:data <=32'hFF2BFFAA;14'd3454:data <=32'hFF0CFFC7;14'd3455:data <=32'hFEF1FFEF;
14'd3456:data <=32'hFF630089;14'd3457:data <=32'hFF6F009B;14'd3458:data <=32'hFF750092;
14'd3459:data <=32'hFF010046;14'd3460:data <=32'hFEC50083;14'd3461:data <=32'hFEDC00C0;
14'd3462:data <=32'hFF0300F9;14'd3463:data <=32'hFF350127;14'd3464:data <=32'hFF73014A;
14'd3465:data <=32'hFFBB015E;14'd3466:data <=32'h0006015F;14'd3467:data <=32'h004E014A;
14'd3468:data <=32'h008B0122;14'd3469:data <=32'h00B800EE;14'd3470:data <=32'h00D300B4;
14'd3471:data <=32'h00D9007A;14'd3472:data <=32'h00D30047;14'd3473:data <=32'h00C2001D;
14'd3474:data <=32'h00AAFFFE;14'd3475:data <=32'h0093FFE8;14'd3476:data <=32'h0078FFDA;
14'd3477:data <=32'h0062FFD2;14'd3478:data <=32'h004AFFCF;14'd3479:data <=32'h0034FFD1;
14'd3480:data <=32'h0021FFD9;14'd3481:data <=32'h0013FFE6;14'd3482:data <=32'h000BFFF6;
14'd3483:data <=32'h000B0007;14'd3484:data <=32'h00110014;14'd3485:data <=32'h001A001C;
14'd3486:data <=32'h0025001F;14'd3487:data <=32'h002E001F;14'd3488:data <=32'h0035001D;
14'd3489:data <=32'h0039001A;14'd3490:data <=32'h003D001A;14'd3491:data <=32'h0045001B;
14'd3492:data <=32'h0050001C;14'd3493:data <=32'h005E0019;14'd3494:data <=32'h006D000F;
14'd3495:data <=32'h007C0000;14'd3496:data <=32'h0088FFEA;14'd3497:data <=32'h008AFFD0;
14'd3498:data <=32'h0086FFB3;14'd3499:data <=32'h0078FF9A;14'd3500:data <=32'h0065FF86;
14'd3501:data <=32'h004DFF79;14'd3502:data <=32'h0036FF73;14'd3503:data <=32'h001FFF73;
14'd3504:data <=32'h000BFF76;14'd3505:data <=32'hFFFBFF7F;14'd3506:data <=32'hFFEDFF89;
14'd3507:data <=32'hFFE2FF95;14'd3508:data <=32'hFFDDFFA3;14'd3509:data <=32'hFFDDFFB0;
14'd3510:data <=32'hFFE4FFBC;14'd3511:data <=32'hFFF1FFC1;14'd3512:data <=32'h0000FFBD;
14'd3513:data <=32'h000EFFAD;14'd3514:data <=32'h0012FF94;14'd3515:data <=32'h000CFF75;
14'd3516:data <=32'hFFF7FF56;14'd3517:data <=32'hFFD2FF3D;14'd3518:data <=32'hFFA3FF2F;
14'd3519:data <=32'hFF6FFF32;14'd3520:data <=32'hFF60FF94;14'd3521:data <=32'hFF3DFF9F;
14'd3522:data <=32'hFF36FFAA;14'd3523:data <=32'hFF59FF83;14'd3524:data <=32'hFEFAFFA6;
14'd3525:data <=32'hFEE9FFD4;14'd3526:data <=32'hFEE20006;14'd3527:data <=32'hFEE50037;
14'd3528:data <=32'hFEF3006B;14'd3529:data <=32'hFF0F0099;14'd3530:data <=32'hFF3500BF;
14'd3531:data <=32'hFF6200D9;14'd3532:data <=32'hFF9100E5;14'd3533:data <=32'hFFBD00E2;
14'd3534:data <=32'hFFE300D9;14'd3535:data <=32'hFFFF00C9;14'd3536:data <=32'h001400B9;
14'd3537:data <=32'h002400AC;14'd3538:data <=32'h003200A1;14'd3539:data <=32'h00410095;
14'd3540:data <=32'h00520089;14'd3541:data <=32'h00610077;14'd3542:data <=32'h006C0062;
14'd3543:data <=32'h0072004B;14'd3544:data <=32'h00720033;14'd3545:data <=32'h006C001D;
14'd3546:data <=32'h0061000B;14'd3547:data <=32'h0054FFFD;14'd3548:data <=32'h0046FFF4;
14'd3549:data <=32'h0038FFED;14'd3550:data <=32'h0028FFEA;14'd3551:data <=32'h0018FFEB;
14'd3552:data <=32'h0005FFF1;14'd3553:data <=32'hFFF5FFFE;14'd3554:data <=32'hFFE90012;
14'd3555:data <=32'hFFE6002B;14'd3556:data <=32'hFFEC0047;14'd3557:data <=32'hFFFD0061;
14'd3558:data <=32'h00190075;14'd3559:data <=32'h003D007E;14'd3560:data <=32'h0063007A;
14'd3561:data <=32'h00860069;14'd3562:data <=32'h00A3004D;14'd3563:data <=32'h00B6002B;
14'd3564:data <=32'h00BD0007;14'd3565:data <=32'h00BBFFE3;14'd3566:data <=32'h00B2FFC5;
14'd3567:data <=32'h00A3FFAA;14'd3568:data <=32'h0090FF94;14'd3569:data <=32'h007AFF84;
14'd3570:data <=32'h0063FF79;14'd3571:data <=32'h004CFF74;14'd3572:data <=32'h0036FF75;
14'd3573:data <=32'h0023FF7B;14'd3574:data <=32'h0016FF84;14'd3575:data <=32'h0011FF91;
14'd3576:data <=32'h0013FF98;14'd3577:data <=32'h001AFF99;14'd3578:data <=32'h0020FF90;
14'd3579:data <=32'h0023FF80;14'd3580:data <=32'h001DFF6B;14'd3581:data <=32'h000BFF55;
14'd3582:data <=32'hFFF0FF43;14'd3583:data <=32'hFFCEFF3B;14'd3584:data <=32'h003CFF58;
14'd3585:data <=32'h001AFF29;14'd3586:data <=32'hFFEEFF1D;14'd3587:data <=32'hFFA7FF7F;
14'd3588:data <=32'hFF56FF93;14'd3589:data <=32'hFF52FFAE;14'd3590:data <=32'hFF51FFC7;
14'd3591:data <=32'hFF54FFDD;14'd3592:data <=32'hFF58FFF2;14'd3593:data <=32'hFF600005;
14'd3594:data <=32'hFF6C0014;14'd3595:data <=32'hFF790020;14'd3596:data <=32'hFF870025;
14'd3597:data <=32'hFF8D0023;14'd3598:data <=32'hFF900021;14'd3599:data <=32'hFF8B0022;
14'd3600:data <=32'hFF820028;14'd3601:data <=32'hFF780037;14'd3602:data <=32'hFF72004F;
14'd3603:data <=32'hFF77006C;14'd3604:data <=32'hFF860089;14'd3605:data <=32'hFFA000A1;
14'd3606:data <=32'hFFC100B2;14'd3607:data <=32'hFFE300B8;14'd3608:data <=32'h000600B2;
14'd3609:data <=32'h002600A6;14'd3610:data <=32'h003F0093;14'd3611:data <=32'h0054007C;
14'd3612:data <=32'h00610061;14'd3613:data <=32'h00680045;14'd3614:data <=32'h00670028;
14'd3615:data <=32'h005C000A;14'd3616:data <=32'h004AFFF3;14'd3617:data <=32'h0030FFE2;
14'd3618:data <=32'h0012FFDE;14'd3619:data <=32'hFFF3FFE4;14'd3620:data <=32'hFFDAFFF7;
14'd3621:data <=32'hFFCA0012;14'd3622:data <=32'hFFC50031;14'd3623:data <=32'hFFCD0051;
14'd3624:data <=32'hFFDF0069;14'd3625:data <=32'hFFF6007B;14'd3626:data <=32'h00110085;
14'd3627:data <=32'h002B0087;14'd3628:data <=32'h00440084;14'd3629:data <=32'h0059007D;
14'd3630:data <=32'h006E0074;14'd3631:data <=32'h00810069;14'd3632:data <=32'h0094005B;
14'd3633:data <=32'h00A6004B;14'd3634:data <=32'h00B60035;14'd3635:data <=32'h00C2001C;
14'd3636:data <=32'h00C90001;14'd3637:data <=32'h00CCFFE5;14'd3638:data <=32'h00CBFFCA;
14'd3639:data <=32'h00C7FFAF;14'd3640:data <=32'h00C1FF95;14'd3641:data <=32'h00B9FF7A;
14'd3642:data <=32'h00ADFF5C;14'd3643:data <=32'h009AFF3C;14'd3644:data <=32'h007EFF1D;
14'd3645:data <=32'h0057FF02;14'd3646:data <=32'h0028FEF1;14'd3647:data <=32'hFFF4FEEF;
14'd3648:data <=32'h0080FFCB;14'd3649:data <=32'h008BFF96;14'd3650:data <=32'h0075FF59;
14'd3651:data <=32'hFFB8FF23;14'd3652:data <=32'hFF59FF45;14'd3653:data <=32'hFF4CFF72;
14'd3654:data <=32'hFF4BFF9C;14'd3655:data <=32'hFF54FFC2;14'd3656:data <=32'hFF63FFDF;
14'd3657:data <=32'hFF76FFF7;14'd3658:data <=32'hFF8E0006;14'd3659:data <=32'hFFA6000D;
14'd3660:data <=32'hFFBE0008;14'd3661:data <=32'hFFD0FFFC;14'd3662:data <=32'hFFD6FFE7;
14'd3663:data <=32'hFFD1FFD3;14'd3664:data <=32'hFFBFFFC2;14'd3665:data <=32'hFFA7FFBB;
14'd3666:data <=32'hFF8BFFC3;14'd3667:data <=32'hFF72FFD5;14'd3668:data <=32'hFF61FFF0;
14'd3669:data <=32'hFF5A0010;14'd3670:data <=32'hFF5F0031;14'd3671:data <=32'hFF6B004C;
14'd3672:data <=32'hFF7E0063;14'd3673:data <=32'hFF940074;14'd3674:data <=32'hFFAB007F;
14'd3675:data <=32'hFFC30085;14'd3676:data <=32'hFFDC0086;14'd3677:data <=32'hFFF30081;
14'd3678:data <=32'h00090078;14'd3679:data <=32'h001B0068;14'd3680:data <=32'h00280055;
14'd3681:data <=32'h002C003F;14'd3682:data <=32'h0028002B;14'd3683:data <=32'h001E001B;
14'd3684:data <=32'h00110012;14'd3685:data <=32'h0003000F;14'd3686:data <=32'hFFF70012;
14'd3687:data <=32'hFFEE0019;14'd3688:data <=32'hFFEA0020;14'd3689:data <=32'hFFE60025;
14'd3690:data <=32'hFFE3002A;14'd3691:data <=32'hFFDE002F;14'd3692:data <=32'hFFD80038;
14'd3693:data <=32'hFFD00046;14'd3694:data <=32'hFFCD0059;14'd3695:data <=32'hFFCE0073;
14'd3696:data <=32'hFFD9008F;14'd3697:data <=32'hFFEE00AA;14'd3698:data <=32'h000E00C0;
14'd3699:data <=32'h003500CE;14'd3700:data <=32'h006000D4;14'd3701:data <=32'h008D00CF;
14'd3702:data <=32'h00BA00BF;14'd3703:data <=32'h00E700A5;14'd3704:data <=32'h010E0082;
14'd3705:data <=32'h01310053;14'd3706:data <=32'h014B001A;14'd3707:data <=32'h0157FFD9;
14'd3708:data <=32'h0153FF92;14'd3709:data <=32'h013CFF4B;14'd3710:data <=32'h0111FF0D;
14'd3711:data <=32'h00D3FEDC;14'd3712:data <=32'h0084FFC5;14'd3713:data <=32'h0094FFA3;
14'd3714:data <=32'h00A7FF72;14'd3715:data <=32'h0093FEEA;14'd3716:data <=32'h0019FEE7;
14'd3717:data <=32'hFFEDFEFB;14'd3718:data <=32'hFFC9FF15;14'd3719:data <=32'hFFB0FF30;
14'd3720:data <=32'hFF9CFF4F;14'd3721:data <=32'hFF90FF6C;14'd3722:data <=32'hFF8BFF8B;
14'd3723:data <=32'hFF8EFFA5;14'd3724:data <=32'hFF98FFBA;14'd3725:data <=32'hFFA4FFC5;
14'd3726:data <=32'hFFB0FFCA;14'd3727:data <=32'hFFB7FFC8;14'd3728:data <=32'hFFB7FFC3;
14'd3729:data <=32'hFFB0FFC1;14'd3730:data <=32'hFFA4FFC3;14'd3731:data <=32'hFF99FFCC;
14'd3732:data <=32'hFF92FFDB;14'd3733:data <=32'hFF90FFEC;14'd3734:data <=32'hFF94FFFB;
14'd3735:data <=32'hFF9D0008;14'd3736:data <=32'hFFA6000E;14'd3737:data <=32'hFFAE0011;
14'd3738:data <=32'hFFB40011;14'd3739:data <=32'hFFB50012;14'd3740:data <=32'hFFB60013;
14'd3741:data <=32'hFFB50017;14'd3742:data <=32'hFFB7001C;14'd3743:data <=32'hFFB90021;
14'd3744:data <=32'hFFBC0026;14'd3745:data <=32'hFFC00028;14'd3746:data <=32'hFFC2002D;
14'd3747:data <=32'hFFC30031;14'd3748:data <=32'hFFC50037;14'd3749:data <=32'hFFCA003E;
14'd3750:data <=32'hFFD20044;14'd3751:data <=32'hFFDF0049;14'd3752:data <=32'hFFEB0048;
14'd3753:data <=32'hFFF80041;14'd3754:data <=32'hFFFF0034;14'd3755:data <=32'h00010024;
14'd3756:data <=32'hFFF80013;14'd3757:data <=32'hFFE60008;14'd3758:data <=32'hFFCE0006;
14'd3759:data <=32'hFFB50010;14'd3760:data <=32'hFF9F0024;14'd3761:data <=32'hFF910043;
14'd3762:data <=32'hFF8C0069;14'd3763:data <=32'hFF950090;14'd3764:data <=32'hFFA800B5;
14'd3765:data <=32'hFFC500D6;14'd3766:data <=32'hFFEC00F1;14'd3767:data <=32'h001A0103;
14'd3768:data <=32'h004D010C;14'd3769:data <=32'h00860109;14'd3770:data <=32'h00C000F6;
14'd3771:data <=32'h00F700D5;14'd3772:data <=32'h012500A3;14'd3773:data <=32'h01450065;
14'd3774:data <=32'h01520021;14'd3775:data <=32'h014DFFDE;14'd3776:data <=32'h010A000C;
14'd3777:data <=32'h011EFFDA;14'd3778:data <=32'h0129FFBA;14'd3779:data <=32'h012BFFD3;
14'd3780:data <=32'h00D9FFAC;14'd3781:data <=32'h00CBFF96;14'd3782:data <=32'h00BDFF82;
14'd3783:data <=32'h00AEFF6D;14'd3784:data <=32'h009AFF56;14'd3785:data <=32'h0081FF43;
14'd3786:data <=32'h0064FF36;14'd3787:data <=32'h0047FF2C;14'd3788:data <=32'h0029FF29;
14'd3789:data <=32'h000CFF29;14'd3790:data <=32'hFFF1FF2B;14'd3791:data <=32'hFFD3FF31;
14'd3792:data <=32'hFFB5FF3B;14'd3793:data <=32'hFF97FF4B;14'd3794:data <=32'hFF7BFF65;
14'd3795:data <=32'hFF64FF87;14'd3796:data <=32'hFF58FFAE;14'd3797:data <=32'hFF5AFFD8;
14'd3798:data <=32'hFF68FFFD;14'd3799:data <=32'hFF82001B;14'd3800:data <=32'hFFA0002B;
14'd3801:data <=32'hFFBF0030;14'd3802:data <=32'hFFDB0029;14'd3803:data <=32'hFFEE001B;
14'd3804:data <=32'hFFFA000A;14'd3805:data <=32'hFFFFFFF8;14'd3806:data <=32'hFFFEFFE7;
14'd3807:data <=32'hFFF6FFD8;14'd3808:data <=32'hFFECFFCC;14'd3809:data <=32'hFFDDFFC4;
14'd3810:data <=32'hFFCCFFBF;14'd3811:data <=32'hFFB8FFC2;14'd3812:data <=32'hFFA5FFCB;
14'd3813:data <=32'hFF96FFDA;14'd3814:data <=32'hFF8CFFEE;14'd3815:data <=32'hFF8A0004;
14'd3816:data <=32'hFF8F0019;14'd3817:data <=32'hFF9B0028;14'd3818:data <=32'hFFA90030;
14'd3819:data <=32'hFFB70030;14'd3820:data <=32'hFFBF002B;14'd3821:data <=32'hFFC10023;
14'd3822:data <=32'hFFBC001D;14'd3823:data <=32'hFFB1001D;14'd3824:data <=32'hFFA40024;
14'd3825:data <=32'hFF990033;14'd3826:data <=32'hFF920045;14'd3827:data <=32'hFF93005B;
14'd3828:data <=32'hFF980071;14'd3829:data <=32'hFFA30087;14'd3830:data <=32'hFFB1009A;
14'd3831:data <=32'hFFC400AC;14'd3832:data <=32'hFFDA00BC;14'd3833:data <=32'hFFF500C8;
14'd3834:data <=32'h001200D0;14'd3835:data <=32'h003500D1;14'd3836:data <=32'h005600C9;
14'd3837:data <=32'h007600B9;14'd3838:data <=32'h009000A1;14'd3839:data <=32'h00A10088;
14'd3840:data <=32'h00D700F5;14'd3841:data <=32'h011200D3;14'd3842:data <=32'h012800A6;
14'd3843:data <=32'h0099008A;14'd3844:data <=32'h0066007F;14'd3845:data <=32'h00800084;
14'd3846:data <=32'h00A00080;14'd3847:data <=32'h00C50073;14'd3848:data <=32'h00E40056;
14'd3849:data <=32'h00FC002F;14'd3850:data <=32'h010A0002;14'd3851:data <=32'h010FFFD2;
14'd3852:data <=32'h0108FFA1;14'd3853:data <=32'h00F7FF72;14'd3854:data <=32'h00DDFF46;
14'd3855:data <=32'h00B7FF20;14'd3856:data <=32'h0088FF00;14'd3857:data <=32'h0050FEEC;
14'd3858:data <=32'h0014FEE7;14'd3859:data <=32'hFFD8FEF5;14'd3860:data <=32'hFFA2FF12;
14'd3861:data <=32'hFF7AFF3E;14'd3862:data <=32'hFF63FF71;14'd3863:data <=32'hFF5DFFA5;
14'd3864:data <=32'hFF67FFD3;14'd3865:data <=32'hFF7BFFF7;14'd3866:data <=32'hFF960010;
14'd3867:data <=32'hFFB1001F;14'd3868:data <=32'hFFCD0024;14'd3869:data <=32'hFFE60023;
14'd3870:data <=32'hFFFC001B;14'd3871:data <=32'h000D0011;14'd3872:data <=32'h001B0001;
14'd3873:data <=32'h0023FFED;14'd3874:data <=32'h0027FFD8;14'd3875:data <=32'h0023FFC1;
14'd3876:data <=32'h0016FFAE;14'd3877:data <=32'h0006FF9E;14'd3878:data <=32'hFFF1FF96;
14'd3879:data <=32'hFFDBFF93;14'd3880:data <=32'hFFC9FF95;14'd3881:data <=32'hFFB8FF99;
14'd3882:data <=32'hFFAAFF9F;14'd3883:data <=32'hFF9BFFA4;14'd3884:data <=32'hFF8CFFAA;
14'd3885:data <=32'hFF78FFB2;14'd3886:data <=32'hFF64FFBE;14'd3887:data <=32'hFF4FFFD2;
14'd3888:data <=32'hFF3DFFEE;14'd3889:data <=32'hFF310011;14'd3890:data <=32'hFF300037;
14'd3891:data <=32'hFF3A005E;14'd3892:data <=32'hFF4F0081;14'd3893:data <=32'hFF6A009C;
14'd3894:data <=32'hFF8900AE;14'd3895:data <=32'hFFA900B9;14'd3896:data <=32'hFFC900BC;
14'd3897:data <=32'hFFE500B9;14'd3898:data <=32'h000000B1;14'd3899:data <=32'h001500A6;
14'd3900:data <=32'h00280095;14'd3901:data <=32'h00340082;14'd3902:data <=32'h0039006D;
14'd3903:data <=32'h0035005C;14'd3904:data <=32'hFFE70104;14'd3905:data <=32'h00170117;
14'd3906:data <=32'h004C0106;14'd3907:data <=32'h0031006C;14'd3908:data <=32'hFFE9006E;
14'd3909:data <=32'hFFF1008B;14'd3910:data <=32'h000500A4;14'd3911:data <=32'h002500B9;
14'd3912:data <=32'h004D00C1;14'd3913:data <=32'h007600BC;14'd3914:data <=32'h009E00AB;
14'd3915:data <=32'h00C10092;14'd3916:data <=32'h00DD0072;14'd3917:data <=32'h00F3004C;
14'd3918:data <=32'h0103001F;14'd3919:data <=32'h0106FFEF;14'd3920:data <=32'h00FEFFBE;
14'd3921:data <=32'h00EAFF8F;14'd3922:data <=32'h00C9FF66;14'd3923:data <=32'h009FFF48;
14'd3924:data <=32'h006FFF39;14'd3925:data <=32'h0041FF38;14'd3926:data <=32'h0019FF43;
14'd3927:data <=32'hFFF8FF58;14'd3928:data <=32'hFFE2FF6E;14'd3929:data <=32'hFFD4FF85;
14'd3930:data <=32'hFFCEFF9A;14'd3931:data <=32'hFFC9FFAB;14'd3932:data <=32'hFFC6FFBC;
14'd3933:data <=32'hFFC5FFCC;14'd3934:data <=32'hFFC6FFDD;14'd3935:data <=32'hFFCDFFEE;
14'd3936:data <=32'hFFD8FFFE;14'd3937:data <=32'hFFE80009;14'd3938:data <=32'hFFFC000F;
14'd3939:data <=32'h0010000D;14'd3940:data <=32'h00230006;14'd3941:data <=32'h0033FFF9;
14'd3942:data <=32'h003FFFE9;14'd3943:data <=32'h0048FFD3;14'd3944:data <=32'h004BFFBD;
14'd3945:data <=32'h004BFFA5;14'd3946:data <=32'h0043FF89;14'd3947:data <=32'h0036FF6C;
14'd3948:data <=32'h001FFF4F;14'd3949:data <=32'hFFFCFF36;14'd3950:data <=32'hFFD1FF25;
14'd3951:data <=32'hFF9EFF22;14'd3952:data <=32'hFF67FF2E;14'd3953:data <=32'hFF35FF4A;
14'd3954:data <=32'hFF0CFF75;14'd3955:data <=32'hFEF0FFA9;14'd3956:data <=32'hFEE4FFE3;
14'd3957:data <=32'hFEE8001B;14'd3958:data <=32'hFEFA004D;14'd3959:data <=32'hFF140077;
14'd3960:data <=32'hFF350098;14'd3961:data <=32'hFF5A00AF;14'd3962:data <=32'hFF8000BC;
14'd3963:data <=32'hFFA700C2;14'd3964:data <=32'hFFCB00BE;14'd3965:data <=32'hFFEB00B0;
14'd3966:data <=32'h0002009D;14'd3967:data <=32'h00100085;14'd3968:data <=32'hFFB60071;
14'd3969:data <=32'hFFB70082;14'd3970:data <=32'hFFCC009A;14'd3971:data <=32'h0013009F;
14'd3972:data <=32'hFFD60090;14'd3973:data <=32'hFFDD009E;14'd3974:data <=32'hFFEF00AC;
14'd3975:data <=32'h000600B8;14'd3976:data <=32'h002400B9;14'd3977:data <=32'h004100B3;
14'd3978:data <=32'h005A00A6;14'd3979:data <=32'h006F0094;14'd3980:data <=32'h007E0080;
14'd3981:data <=32'h0089006C;14'd3982:data <=32'h00930058;14'd3983:data <=32'h00990043;
14'd3984:data <=32'h009D002C;14'd3985:data <=32'h009B0016;14'd3986:data <=32'h0095FFFF;
14'd3987:data <=32'h0089FFEE;14'd3988:data <=32'h007AFFE0;14'd3989:data <=32'h006BFFDB;
14'd3990:data <=32'h0061FFD9;14'd3991:data <=32'h005AFFDA;14'd3992:data <=32'h0058FFDA;
14'd3993:data <=32'h005AFFD7;14'd3994:data <=32'h005CFFCD;14'd3995:data <=32'h0059FFC0;
14'd3996:data <=32'h0050FFB1;14'd3997:data <=32'h0041FFA5;14'd3998:data <=32'h002DFF9E;
14'd3999:data <=32'h0016FF9F;14'd4000:data <=32'h0003FFA8;14'd4001:data <=32'hFFF3FFB7;
14'd4002:data <=32'hFFEAFFC9;14'd4003:data <=32'hFFE9FFDD;14'd4004:data <=32'hFFEFFFEF;
14'd4005:data <=32'hFFF8FFFE;14'd4006:data <=32'h00080008;14'd4007:data <=32'h001C000F;
14'd4008:data <=32'h00300010;14'd4009:data <=32'h00490009;14'd4010:data <=32'h0061FFF9;
14'd4011:data <=32'h0075FFE0;14'd4012:data <=32'h0082FFBD;14'd4013:data <=32'h0084FF94;
14'd4014:data <=32'h0078FF69;14'd4015:data <=32'h005EFF40;14'd4016:data <=32'h0036FF21;
14'd4017:data <=32'h0005FF0F;14'd4018:data <=32'hFFD3FF0B;14'd4019:data <=32'hFFA3FF15;
14'd4020:data <=32'hFF78FF2A;14'd4021:data <=32'hFF57FF47;14'd4022:data <=32'hFF3EFF67;
14'd4023:data <=32'hFF2CFF87;14'd4024:data <=32'hFF20FFA8;14'd4025:data <=32'hFF19FFC9;
14'd4026:data <=32'hFF17FFE9;14'd4027:data <=32'hFF19000A;14'd4028:data <=32'hFF200029;
14'd4029:data <=32'hFF2D0043;14'd4030:data <=32'hFF3E005B;14'd4031:data <=32'hFF4E006B;
14'd4032:data <=32'hFFC4006D;14'd4033:data <=32'hFFC80061;14'd4034:data <=32'hFFB70063;
14'd4035:data <=32'hFF4B00A0;14'd4036:data <=32'hFF1C00AF;14'd4037:data <=32'hFF3B00D9;
14'd4038:data <=32'hFF6500FD;14'd4039:data <=32'hFF980117;14'd4040:data <=32'hFFD30121;
14'd4041:data <=32'h000D0119;14'd4042:data <=32'h00410103;14'd4043:data <=32'h006A00E0;
14'd4044:data <=32'h008600B9;14'd4045:data <=32'h00950090;14'd4046:data <=32'h0099006A;
14'd4047:data <=32'h00950046;14'd4048:data <=32'h008C0028;14'd4049:data <=32'h007C000F;
14'd4050:data <=32'h0067FFFC;14'd4051:data <=32'h004FFFF2;14'd4052:data <=32'h0037FFF0;
14'd4053:data <=32'h0022FFF8;14'd4054:data <=32'h00120008;14'd4055:data <=32'h000D001D;
14'd4056:data <=32'h00140031;14'd4057:data <=32'h0024003F;14'd4058:data <=32'h003A0044;
14'd4059:data <=32'h00510040;14'd4060:data <=32'h00630031;14'd4061:data <=32'h006E001E;
14'd4062:data <=32'h00710008;14'd4063:data <=32'h006DFFF4;14'd4064:data <=32'h0062FFE5;
14'd4065:data <=32'h0056FFDB;14'd4066:data <=32'h004AFFD6;14'd4067:data <=32'h003EFFD5;
14'd4068:data <=32'h0036FFD6;14'd4069:data <=32'h002FFFD9;14'd4070:data <=32'h002AFFDE;
14'd4071:data <=32'h0026FFE4;14'd4072:data <=32'h0027FFEB;14'd4073:data <=32'h002BFFF2;
14'd4074:data <=32'h0035FFF8;14'd4075:data <=32'h0043FFF8;14'd4076:data <=32'h0051FFF2;
14'd4077:data <=32'h005EFFE5;14'd4078:data <=32'h0067FFD3;14'd4079:data <=32'h006AFFBC;
14'd4080:data <=32'h0065FFA5;14'd4081:data <=32'h005AFF92;14'd4082:data <=32'h004BFF84;
14'd4083:data <=32'h003CFF7B;14'd4084:data <=32'h002FFF74;14'd4085:data <=32'h0024FF6E;
14'd4086:data <=32'h001DFF68;14'd4087:data <=32'h0012FF5B;14'd4088:data <=32'h0004FF4C;
14'd4089:data <=32'hFFEFFF3D;14'd4090:data <=32'hFFD3FF30;14'd4091:data <=32'hFFB0FF2A;
14'd4092:data <=32'hFF8BFF2B;14'd4093:data <=32'hFF63FF35;14'd4094:data <=32'hFF3DFF47;
14'd4095:data <=32'hFF19FF60;14'd4096:data <=32'hFF630020;14'd4097:data <=32'hFF670022;
14'd4098:data <=32'hFF63000C;14'd4099:data <=32'hFEF3FF9C;14'd4100:data <=32'hFE97FFC0;
14'd4101:data <=32'hFE8C000B;14'd4102:data <=32'hFE950059;14'd4103:data <=32'hFEB200A3;
14'd4104:data <=32'hFEE300E0;14'd4105:data <=32'hFF23010C;14'd4106:data <=32'hFF680123;
14'd4107:data <=32'hFFAA0127;14'd4108:data <=32'hFFE7011B;14'd4109:data <=32'h00180104;
14'd4110:data <=32'h004100E5;14'd4111:data <=32'h005E00C1;14'd4112:data <=32'h0071009B;
14'd4113:data <=32'h007B0076;14'd4114:data <=32'h007C0050;14'd4115:data <=32'h0072002E;
14'd4116:data <=32'h005F0015;14'd4117:data <=32'h00470003;14'd4118:data <=32'h002EFFFD;
14'd4119:data <=32'h00170002;14'd4120:data <=32'h0008000E;14'd4121:data <=32'h0002001D;
14'd4122:data <=32'h0002002B;14'd4123:data <=32'h000A0034;14'd4124:data <=32'h00130039;
14'd4125:data <=32'h001A0039;14'd4126:data <=32'h001F0037;14'd4127:data <=32'h00210037;
14'd4128:data <=32'h00220038;14'd4129:data <=32'h0026003C;14'd4130:data <=32'h002B0040;
14'd4131:data <=32'h00360044;14'd4132:data <=32'h00430045;14'd4133:data <=32'h00520041;
14'd4134:data <=32'h005E0039;14'd4135:data <=32'h006A002C;14'd4136:data <=32'h0070001E;
14'd4137:data <=32'h00750011;14'd4138:data <=32'h00770002;14'd4139:data <=32'h0078FFF4;
14'd4140:data <=32'h0077FFE6;14'd4141:data <=32'h0073FFD7;14'd4142:data <=32'h006CFFC9;
14'd4143:data <=32'h0060FFBB;14'd4144:data <=32'h0051FFB3;14'd4145:data <=32'h0040FFB0;
14'd4146:data <=32'h0032FFB6;14'd4147:data <=32'h0027FFC1;14'd4148:data <=32'h0026FFCE;
14'd4149:data <=32'h002FFFDB;14'd4150:data <=32'h0041FFE2;14'd4151:data <=32'h0057FFDD;
14'd4152:data <=32'h006DFFCD;14'd4153:data <=32'h007FFFB0;14'd4154:data <=32'h0085FF8C;
14'd4155:data <=32'h007FFF63;14'd4156:data <=32'h006EFF3B;14'd4157:data <=32'h0050FF17;
14'd4158:data <=32'h0028FEF9;14'd4159:data <=32'hFFF8FEE4;14'd4160:data <=32'hFFBEFF59;
14'd4161:data <=32'hFFA5FF47;14'd4162:data <=32'hFF9DFF3D;14'd4163:data <=32'hFFBFFF03;
14'd4164:data <=32'hFF48FEFA;14'd4165:data <=32'hFF15FF20;14'd4166:data <=32'hFEEEFF55;
14'd4167:data <=32'hFED5FF91;14'd4168:data <=32'hFECFFFCF;14'd4169:data <=32'hFEDB0007;
14'd4170:data <=32'hFEF10037;14'd4171:data <=32'hFF0D005B;14'd4172:data <=32'hFF2C0077;
14'd4173:data <=32'hFF4A0089;14'd4174:data <=32'hFF660098;14'd4175:data <=32'hFF8200A2;
14'd4176:data <=32'hFF9F00A8;14'd4177:data <=32'hFFBB00AA;14'd4178:data <=32'hFFD800A7;
14'd4179:data <=32'hFFF1009E;14'd4180:data <=32'h00060090;14'd4181:data <=32'h00150082;
14'd4182:data <=32'h001E0071;14'd4183:data <=32'h00240065;14'd4184:data <=32'h002A0059;
14'd4185:data <=32'h002F004E;14'd4186:data <=32'h00350042;14'd4187:data <=32'h00380032;
14'd4188:data <=32'h00370021;14'd4189:data <=32'h00300010;14'd4190:data <=32'h00200001;
14'd4191:data <=32'h000CFFF9;14'd4192:data <=32'hFFF5FFFA;14'd4193:data <=32'hFFDF0007;
14'd4194:data <=32'hFFCF001A;14'd4195:data <=32'hFFC80035;14'd4196:data <=32'hFFCB0051;
14'd4197:data <=32'hFFD80069;14'd4198:data <=32'hFFEE007F;14'd4199:data <=32'h0007008B;
14'd4200:data <=32'h00240090;14'd4201:data <=32'h0040008E;14'd4202:data <=32'h005B0086;
14'd4203:data <=32'h00760079;14'd4204:data <=32'h008B0063;14'd4205:data <=32'h009C004A;
14'd4206:data <=32'h00A7002E;14'd4207:data <=32'h00A8000F;14'd4208:data <=32'h00A0FFF2;
14'd4209:data <=32'h008FFFDA;14'd4210:data <=32'h007BFFCC;14'd4211:data <=32'h0065FFC7;
14'd4212:data <=32'h0054FFCC;14'd4213:data <=32'h004AFFD8;14'd4214:data <=32'h004CFFE3;
14'd4215:data <=32'h0056FFEC;14'd4216:data <=32'h0066FFEC;14'd4217:data <=32'h007AFFE3;
14'd4218:data <=32'h0088FFD0;14'd4219:data <=32'h0092FFB6;14'd4220:data <=32'h0092FF99;
14'd4221:data <=32'h008CFF7B;14'd4222:data <=32'h007FFF5F;14'd4223:data <=32'h006BFF44;
14'd4224:data <=32'h00AAFF87;14'd4225:data <=32'h00AAFF47;14'd4226:data <=32'h0090FF1E;
14'd4227:data <=32'h003BFF50;14'd4228:data <=32'hFFDEFF30;14'd4229:data <=32'hFFC0FF3C;
14'd4230:data <=32'hFFA7FF4F;14'd4231:data <=32'hFF93FF66;14'd4232:data <=32'hFF89FF7E;
14'd4233:data <=32'hFF88FF94;14'd4234:data <=32'hFF8AFFA2;14'd4235:data <=32'hFF8DFFAA;
14'd4236:data <=32'hFF8BFFAD;14'd4237:data <=32'hFF83FFAD;14'd4238:data <=32'hFF75FFB2;
14'd4239:data <=32'hFF64FFBE;14'd4240:data <=32'hFF54FFD0;14'd4241:data <=32'hFF47FFE9;
14'd4242:data <=32'hFF440006;14'd4243:data <=32'hFF450024;14'd4244:data <=32'hFF4E0041;
14'd4245:data <=32'hFF5B005B;14'd4246:data <=32'hFF6F0073;14'd4247:data <=32'hFF850088;
14'd4248:data <=32'hFFA20099;14'd4249:data <=32'hFFC400A2;14'd4250:data <=32'hFFE800A3;
14'd4251:data <=32'h000C0099;14'd4252:data <=32'h002C0082;14'd4253:data <=32'h00420064;
14'd4254:data <=32'h004D0040;14'd4255:data <=32'h0048001B;14'd4256:data <=32'h0037FFFC;
14'd4257:data <=32'h001CFFE7;14'd4258:data <=32'hFFFEFFE0;14'd4259:data <=32'hFFE1FFE3;
14'd4260:data <=32'hFFC7FFF1;14'd4261:data <=32'hFFB50005;14'd4262:data <=32'hFFAA001D;
14'd4263:data <=32'hFFA60036;14'd4264:data <=32'hFFA9004D;14'd4265:data <=32'hFFB10065;
14'd4266:data <=32'hFFBF007B;14'd4267:data <=32'hFFD1008D;14'd4268:data <=32'hFFE7009E;
14'd4269:data <=32'h000200A7;14'd4270:data <=32'h001F00AA;14'd4271:data <=32'h003B00A6;
14'd4272:data <=32'h0054009C;14'd4273:data <=32'h0069008E;14'd4274:data <=32'h0079007F;
14'd4275:data <=32'h00840071;14'd4276:data <=32'h008F0066;14'd4277:data <=32'h009B005B;
14'd4278:data <=32'h00AA0050;14'd4279:data <=32'h00BD0041;14'd4280:data <=32'h00CF002A;
14'd4281:data <=32'h00DF000C;14'd4282:data <=32'h00E7FFE7;14'd4283:data <=32'h00E7FFBE;
14'd4284:data <=32'h00DAFF96;14'd4285:data <=32'h00C4FF73;14'd4286:data <=32'h00A7FF57;
14'd4287:data <=32'h0086FF45;14'd4288:data <=32'h00B20039;14'd4289:data <=32'h00E5000A;
14'd4290:data <=32'h00F7FFC2;14'd4291:data <=32'h005AFF48;14'd4292:data <=32'hFFF9FF30;
14'd4293:data <=32'hFFDAFF48;14'd4294:data <=32'hFFC4FF65;14'd4295:data <=32'hFFB9FF85;
14'd4296:data <=32'hFFBBFFA5;14'd4297:data <=32'hFFC8FFBD;14'd4298:data <=32'hFFDDFFCB;
14'd4299:data <=32'hFFF3FFCC;14'd4300:data <=32'h0004FFBF;14'd4301:data <=32'h000BFFAA;
14'd4302:data <=32'h0007FF92;14'd4303:data <=32'hFFF7FF7E;14'd4304:data <=32'hFFDEFF70;
14'd4305:data <=32'hFFC0FF6B;14'd4306:data <=32'hFFA1FF71;14'd4307:data <=32'hFF86FF7E;
14'd4308:data <=32'hFF6EFF91;14'd4309:data <=32'hFF5BFFAA;14'd4310:data <=32'hFF4CFFC8;
14'd4311:data <=32'hFF44FFE8;14'd4312:data <=32'hFF44000C;14'd4313:data <=32'hFF4E002F;
14'd4314:data <=32'hFF610050;14'd4315:data <=32'hFF7E0068;14'd4316:data <=32'hFFA00077;
14'd4317:data <=32'hFFC40079;14'd4318:data <=32'hFFE3006F;14'd4319:data <=32'hFFFB005E;
14'd4320:data <=32'h00080047;14'd4321:data <=32'h000E0032;14'd4322:data <=32'h000C001F;
14'd4323:data <=32'h00050012;14'd4324:data <=32'hFFFC0009;14'd4325:data <=32'hFFF30003;
14'd4326:data <=32'hFFEAFFFE;14'd4327:data <=32'hFFE1FFFA;14'd4328:data <=32'hFFD5FFF7;
14'd4329:data <=32'hFFC8FFF6;14'd4330:data <=32'hFFB8FFFB;14'd4331:data <=32'hFFA60004;
14'd4332:data <=32'hFF970014;14'd4333:data <=32'hFF8A002A;14'd4334:data <=32'hFF830044;
14'd4335:data <=32'hFF820060;14'd4336:data <=32'hFF88007D;14'd4337:data <=32'hFF930099;
14'd4338:data <=32'hFFA400B6;14'd4339:data <=32'hFFBA00D3;14'd4340:data <=32'hFFD800ED;
14'd4341:data <=32'h00000104;14'd4342:data <=32'h00300115;14'd4343:data <=32'h0069011A;
14'd4344:data <=32'h00A7010E;14'd4345:data <=32'h00E300F1;14'd4346:data <=32'h011700C4;
14'd4347:data <=32'h013D0086;14'd4348:data <=32'h01520043;14'd4349:data <=32'h0153FFFE;
14'd4350:data <=32'h0143FFBD;14'd4351:data <=32'h0125FF85;14'd4352:data <=32'h007D0048;
14'd4353:data <=32'h00AB003D;14'd4354:data <=32'h00E20016;14'd4355:data <=32'h0107FF77;
14'd4356:data <=32'h00A1FF3B;14'd4357:data <=32'h0073FF35;14'd4358:data <=32'h0046FF3B;
14'd4359:data <=32'h0021FF4A;14'd4360:data <=32'h0007FF62;14'd4361:data <=32'hFFF9FF7D;
14'd4362:data <=32'hFFF8FF95;14'd4363:data <=32'hFFFFFFA5;14'd4364:data <=32'h0009FFAB;
14'd4365:data <=32'h0011FFA7;14'd4366:data <=32'h0014FF9E;14'd4367:data <=32'h0010FF93;
14'd4368:data <=32'h0004FF8A;14'd4369:data <=32'hFFF5FF87;14'd4370:data <=32'hFFE6FF86;
14'd4371:data <=32'hFFD8FF8B;14'd4372:data <=32'hFFCCFF92;14'd4373:data <=32'hFFC1FF97;
14'd4374:data <=32'hFFB7FF9F;14'd4375:data <=32'hFFADFFA9;14'd4376:data <=32'hFFA3FFB3;
14'd4377:data <=32'hFF9DFFC2;14'd4378:data <=32'hFF98FFD3;14'd4379:data <=32'hFF9AFFE2;
14'd4380:data <=32'hFF9FFFF0;14'd4381:data <=32'hFFA8FFF9;14'd4382:data <=32'hFFB1FFFE;
14'd4383:data <=32'hFFB6FFFF;14'd4384:data <=32'hFFB90000;14'd4385:data <=32'hFFB70000;
14'd4386:data <=32'hFFB60005;14'd4387:data <=32'hFFB4000D;14'd4388:data <=32'hFFB80018;
14'd4389:data <=32'hFFC00021;14'd4390:data <=32'hFFCC0027;14'd4391:data <=32'hFFDC0026;
14'd4392:data <=32'hFFEA001E;14'd4393:data <=32'hFFF3000F;14'd4394:data <=32'hFFF4FFFE;
14'd4395:data <=32'hFFEDFFEA;14'd4396:data <=32'hFFDEFFDB;14'd4397:data <=32'hFFC8FFD2;
14'd4398:data <=32'hFFB0FFCF;14'd4399:data <=32'hFF94FFD5;14'd4400:data <=32'hFF78FFE2;
14'd4401:data <=32'hFF5FFFF7;14'd4402:data <=32'hFF490015;14'd4403:data <=32'hFF38003C;
14'd4404:data <=32'hFF30006B;14'd4405:data <=32'hFF3400A1;14'd4406:data <=32'hFF4900D7;
14'd4407:data <=32'hFF6F010A;14'd4408:data <=32'hFFA50134;14'd4409:data <=32'hFFE7014C;
14'd4410:data <=32'h002E0152;14'd4411:data <=32'h00740143;14'd4412:data <=32'h00B20123;
14'd4413:data <=32'h00E300F8;14'd4414:data <=32'h010600C3;14'd4415:data <=32'h011B008D;
14'd4416:data <=32'h00B40093;14'd4417:data <=32'h00DD0081;14'd4418:data <=32'h01020077;
14'd4419:data <=32'h01200087;14'd4420:data <=32'h00ED003A;14'd4421:data <=32'h00EB0017;
14'd4422:data <=32'h00E4FFF9;14'd4423:data <=32'h00D9FFDE;14'd4424:data <=32'h00CCFFC8;
14'd4425:data <=32'h00C0FFB6;14'd4426:data <=32'h00B5FFA6;14'd4427:data <=32'h00ACFF95;
14'd4428:data <=32'h00A0FF7E;14'd4429:data <=32'h0090FF68;14'd4430:data <=32'h0077FF53;
14'd4431:data <=32'h0057FF40;14'd4432:data <=32'h0031FF37;14'd4433:data <=32'h000AFF3C;
14'd4434:data <=32'hFFE6FF4A;14'd4435:data <=32'hFFC9FF62;14'd4436:data <=32'hFFB8FF7E;
14'd4437:data <=32'hFFAFFF9A;14'd4438:data <=32'hFFAFFFB4;14'd4439:data <=32'hFFB4FFCB;
14'd4440:data <=32'hFFBEFFDC;14'd4441:data <=32'hFFCAFFE8;14'd4442:data <=32'hFFD8FFF1;
14'd4443:data <=32'hFFE7FFF5;14'd4444:data <=32'hFFF6FFF3;14'd4445:data <=32'h0004FFEA;
14'd4446:data <=32'h000DFFDC;14'd4447:data <=32'h0010FFC9;14'd4448:data <=32'h0009FFB7;
14'd4449:data <=32'hFFFAFFA7;14'd4450:data <=32'hFFE6FF9F;14'd4451:data <=32'hFFCFFFA1;
14'd4452:data <=32'hFFBAFFAA;14'd4453:data <=32'hFFACFFBB;14'd4454:data <=32'hFFA5FFCE;
14'd4455:data <=32'hFFA7FFE0;14'd4456:data <=32'hFFAFFFEE;14'd4457:data <=32'hFFBAFFF4;
14'd4458:data <=32'hFFC4FFF3;14'd4459:data <=32'hFFCAFFEE;14'd4460:data <=32'hFFCCFFE7;
14'd4461:data <=32'hFFC8FFDF;14'd4462:data <=32'hFFC0FFD9;14'd4463:data <=32'hFFB5FFD4;
14'd4464:data <=32'hFFA7FFD2;14'd4465:data <=32'hFF96FFD4;14'd4466:data <=32'hFF83FFDA;
14'd4467:data <=32'hFF6FFFE6;14'd4468:data <=32'hFF5AFFF9;14'd4469:data <=32'hFF480014;
14'd4470:data <=32'hFF3E0037;14'd4471:data <=32'hFF3D0060;14'd4472:data <=32'hFF490088;
14'd4473:data <=32'hFF6100AC;14'd4474:data <=32'hFF8100C8;14'd4475:data <=32'hFFA600D9;
14'd4476:data <=32'hFFCA00E1;14'd4477:data <=32'hFFEA00E0;14'd4478:data <=32'h000600DB;
14'd4479:data <=32'h001D00D6;14'd4480:data <=32'h00310134;14'd4481:data <=32'h006F013A;
14'd4482:data <=32'h00960129;14'd4483:data <=32'h002900F6;14'd4484:data <=32'h000E00D6;
14'd4485:data <=32'h002E00DE;14'd4486:data <=32'h005100E1;14'd4487:data <=32'h007800DB;
14'd4488:data <=32'h009C00D0;14'd4489:data <=32'h00C200BD;14'd4490:data <=32'h00E800A2;
14'd4491:data <=32'h010A007B;14'd4492:data <=32'h0125004B;14'd4493:data <=32'h01330011;
14'd4494:data <=32'h0132FFD0;14'd4495:data <=32'h011DFF92;14'd4496:data <=32'h00F8FF5C;
14'd4497:data <=32'h00C5FF33;14'd4498:data <=32'h008BFF1C;14'd4499:data <=32'h0051FF19;
14'd4500:data <=32'h001CFF24;14'd4501:data <=32'hFFF1FF3A;14'd4502:data <=32'hFFD1FF57;
14'd4503:data <=32'hFFBAFF78;14'd4504:data <=32'hFFADFF9B;14'd4505:data <=32'hFFABFFBC;
14'd4506:data <=32'hFFB0FFDC;14'd4507:data <=32'hFFBDFFF8;14'd4508:data <=32'hFFD3000D;
14'd4509:data <=32'hFFED0019;14'd4510:data <=32'h0009001C;14'd4511:data <=32'h00230013;
14'd4512:data <=32'h00370001;14'd4513:data <=32'h0043FFEC;14'd4514:data <=32'h0045FFD3;
14'd4515:data <=32'h003FFFBE;14'd4516:data <=32'h0034FFAF;14'd4517:data <=32'h0028FFA5;
14'd4518:data <=32'h001AFF9D;14'd4519:data <=32'h0011FF99;14'd4520:data <=32'h0008FF94;
14'd4521:data <=32'h0000FF8D;14'd4522:data <=32'hFFF5FF85;14'd4523:data <=32'hFFE6FF7E;
14'd4524:data <=32'hFFD2FF78;14'd4525:data <=32'hFFBAFF77;14'd4526:data <=32'hFFA3FF7B;
14'd4527:data <=32'hFF8BFF86;14'd4528:data <=32'hFF76FF97;14'd4529:data <=32'hFF67FFAB;
14'd4530:data <=32'hFF5BFFC1;14'd4531:data <=32'hFF53FFD9;14'd4532:data <=32'hFF4EFFF0;
14'd4533:data <=32'hFF4C0008;14'd4534:data <=32'hFF4F0023;14'd4535:data <=32'hFF59003C;
14'd4536:data <=32'hFF680054;14'd4537:data <=32'hFF7D0064;14'd4538:data <=32'hFF96006E;
14'd4539:data <=32'hFFAC006E;14'd4540:data <=32'hFFBE0065;14'd4541:data <=32'hFFC70059;
14'd4542:data <=32'hFFC6004D;14'd4543:data <=32'hFFBB0047;14'd4544:data <=32'hFF4D00CF;
14'd4545:data <=32'hFF6900FF;14'd4546:data <=32'hFF9C010E;14'd4547:data <=32'hFFB1007B;
14'd4548:data <=32'hFF78006A;14'd4549:data <=32'hFF7C008D;14'd4550:data <=32'hFF8900B0;
14'd4551:data <=32'hFFA100D0;14'd4552:data <=32'hFFC100EC;14'd4553:data <=32'hFFE90103;
14'd4554:data <=32'h00180112;14'd4555:data <=32'h00500114;14'd4556:data <=32'h00890107;
14'd4557:data <=32'h00BF00E8;14'd4558:data <=32'h00EC00BC;14'd4559:data <=32'h01090084;
14'd4560:data <=32'h01160047;14'd4561:data <=32'h010F000C;14'd4562:data <=32'h00FCFFD9;
14'd4563:data <=32'h00DEFFB0;14'd4564:data <=32'h00BAFF95;14'd4565:data <=32'h0097FF83;
14'd4566:data <=32'h0076FF7A;14'd4567:data <=32'h0056FF77;14'd4568:data <=32'h0039FF79;
14'd4569:data <=32'h001EFF80;14'd4570:data <=32'h0005FF8E;14'd4571:data <=32'hFFF2FFA0;
14'd4572:data <=32'hFFE4FFB5;14'd4573:data <=32'hFFDFFFCD;14'd4574:data <=32'hFFE1FFE3;
14'd4575:data <=32'hFFE9FFF6;14'd4576:data <=32'hFFF60003;14'd4577:data <=32'h0003000C;
14'd4578:data <=32'h00110011;14'd4579:data <=32'h001D0012;14'd4580:data <=32'h002B0012;
14'd4581:data <=32'h003B0010;14'd4582:data <=32'h004B000D;14'd4583:data <=32'h005F0003;
14'd4584:data <=32'h0072FFF2;14'd4585:data <=32'h0083FFD7;14'd4586:data <=32'h008DFFB4;
14'd4587:data <=32'h008BFF8D;14'd4588:data <=32'h007DFF64;14'd4589:data <=32'h0062FF3F;
14'd4590:data <=32'h003DFF22;14'd4591:data <=32'h000EFF11;14'd4592:data <=32'hFFDEFF0B;
14'd4593:data <=32'hFFAEFF13;14'd4594:data <=32'hFF83FF24;14'd4595:data <=32'hFF5EFF40;
14'd4596:data <=32'hFF3FFF60;14'd4597:data <=32'hFF28FF88;14'd4598:data <=32'hFF1AFFB2;
14'd4599:data <=32'hFF17FFDF;14'd4600:data <=32'hFF21000A;14'd4601:data <=32'hFF360030;
14'd4602:data <=32'hFF53004B;14'd4603:data <=32'hFF75005A;14'd4604:data <=32'hFF96005B;
14'd4605:data <=32'hFFB00050;14'd4606:data <=32'hFFBE003D;14'd4607:data <=32'hFFBF002A;
14'd4608:data <=32'hFF6B000A;14'd4609:data <=32'hFF55001F;14'd4610:data <=32'hFF590046;
14'd4611:data <=32'hFFA40062;14'd4612:data <=32'hFF6E0043;14'd4613:data <=32'hFF700058;
14'd4614:data <=32'hFF76006F;14'd4615:data <=32'hFF820083;14'd4616:data <=32'hFF900096;
14'd4617:data <=32'hFFA300AA;14'd4618:data <=32'hFFB900BA;14'd4619:data <=32'hFFD600C8;
14'd4620:data <=32'hFFF600D0;14'd4621:data <=32'h001A00CD;14'd4622:data <=32'h003C00C1;
14'd4623:data <=32'h005A00AD;14'd4624:data <=32'h006D0093;14'd4625:data <=32'h00770078;
14'd4626:data <=32'h0079005F;14'd4627:data <=32'h0076004D;14'd4628:data <=32'h00730040;
14'd4629:data <=32'h00720037;14'd4630:data <=32'h0073002F;14'd4631:data <=32'h00770025;
14'd4632:data <=32'h007B0018;14'd4633:data <=32'h007D0006;14'd4634:data <=32'h0079FFF4;
14'd4635:data <=32'h0070FFE4;14'd4636:data <=32'h0063FFD7;14'd4637:data <=32'h0054FFCD;
14'd4638:data <=32'h0045FFC7;14'd4639:data <=32'h0036FFC5;14'd4640:data <=32'h0026FFC6;
14'd4641:data <=32'h0017FFCB;14'd4642:data <=32'h0008FFD3;14'd4643:data <=32'hFFFCFFE2;
14'd4644:data <=32'hFFF4FFF4;14'd4645:data <=32'hFFF3000B;14'd4646:data <=32'hFFFC0024;
14'd4647:data <=32'h000F003B;14'd4648:data <=32'h002C004A;14'd4649:data <=32'h0052004E;
14'd4650:data <=32'h00780043;14'd4651:data <=32'h009B002B;14'd4652:data <=32'h00B50006;
14'd4653:data <=32'h00C4FFDB;14'd4654:data <=32'h00C5FFAB;14'd4655:data <=32'h00B8FF7F;
14'd4656:data <=32'h00A0FF57;14'd4657:data <=32'h0081FF37;14'd4658:data <=32'h005DFF20;
14'd4659:data <=32'h0035FF0F;14'd4660:data <=32'h000CFF07;14'd4661:data <=32'hFFE1FF09;
14'd4662:data <=32'hFFB7FF12;14'd4663:data <=32'hFF92FF25;14'd4664:data <=32'hFF73FF3F;
14'd4665:data <=32'hFF5EFF5F;14'd4666:data <=32'hFF51FF80;14'd4667:data <=32'hFF4EFF9D;
14'd4668:data <=32'hFF52FFB5;14'd4669:data <=32'hFF55FFC5;14'd4670:data <=32'hFF57FFD0;
14'd4671:data <=32'hFF54FFD9;14'd4672:data <=32'hFFBB0005;14'd4673:data <=32'hFFB3FFF2;
14'd4674:data <=32'hFF95FFF0;14'd4675:data <=32'hFF1F0017;14'd4676:data <=32'hFEED0015;
14'd4677:data <=32'hFEF70046;14'd4678:data <=32'hFF0E0071;14'd4679:data <=32'hFF2D0095;
14'd4680:data <=32'hFF5300AE;14'd4681:data <=32'hFF7800BF;14'd4682:data <=32'hFF9E00C8;
14'd4683:data <=32'hFFC400C9;14'd4684:data <=32'hFFE800C3;14'd4685:data <=32'h000900B5;
14'd4686:data <=32'h0026009E;14'd4687:data <=32'h00390081;14'd4688:data <=32'h00400062;
14'd4689:data <=32'h003B0045;14'd4690:data <=32'h002D002F;14'd4691:data <=32'h00190024;
14'd4692:data <=32'h00040026;14'd4693:data <=32'hFFF60032;14'd4694:data <=32'hFFF10042;
14'd4695:data <=32'hFFF60055;14'd4696:data <=32'h00030063;14'd4697:data <=32'h0015006B;
14'd4698:data <=32'h0028006B;14'd4699:data <=32'h003B0066;14'd4700:data <=32'h004A005B;
14'd4701:data <=32'h0057004D;14'd4702:data <=32'h005F003E;14'd4703:data <=32'h0064002D;
14'd4704:data <=32'h0066001B;14'd4705:data <=32'h00610009;14'd4706:data <=32'h0057FFF9;
14'd4707:data <=32'h0048FFED;14'd4708:data <=32'h0036FFE8;14'd4709:data <=32'h0024FFEC;
14'd4710:data <=32'h0014FFF7;14'd4711:data <=32'h000C0009;14'd4712:data <=32'h000D001D;
14'd4713:data <=32'h0017002F;14'd4714:data <=32'h002A003D;14'd4715:data <=32'h00400041;
14'd4716:data <=32'h0058003E;14'd4717:data <=32'h006D0033;14'd4718:data <=32'h007C0023;
14'd4719:data <=32'h00870010;14'd4720:data <=32'h008EFFFE;14'd4721:data <=32'h0092FFED;
14'd4722:data <=32'h0095FFDB;14'd4723:data <=32'h0098FFC9;14'd4724:data <=32'h0099FFB3;
14'd4725:data <=32'h0099FF9C;14'd4726:data <=32'h0092FF83;14'd4727:data <=32'h0085FF69;
14'd4728:data <=32'h0075FF51;14'd4729:data <=32'h0062FF3C;14'd4730:data <=32'h004BFF2A;
14'd4731:data <=32'h0032FF1A;14'd4732:data <=32'h0017FF0B;14'd4733:data <=32'hFFF5FEFC;
14'd4734:data <=32'hFFCEFEF1;14'd4735:data <=32'hFF9FFEEC;14'd4736:data <=32'hFF9FFFCA;
14'd4737:data <=32'hFFA0FFBF;14'd4738:data <=32'hFF9BFFA1;14'd4739:data <=32'hFF44FF15;
14'd4740:data <=32'hFEE2FF15;14'd4741:data <=32'hFEBCFF57;14'd4742:data <=32'hFEA9FF9F;
14'd4743:data <=32'hFEAAFFE5;14'd4744:data <=32'hFEBB0027;14'd4745:data <=32'hFED8005E;
14'd4746:data <=32'hFEFD008B;14'd4747:data <=32'hFF2A00AF;14'd4748:data <=32'hFF5D00C6;
14'd4749:data <=32'hFF9100D0;14'd4750:data <=32'hFFC400CC;14'd4751:data <=32'hFFF100BA;
14'd4752:data <=32'h0014009C;14'd4753:data <=32'h00280078;14'd4754:data <=32'h002D0054;
14'd4755:data <=32'h00250035;14'd4756:data <=32'h00160021;14'd4757:data <=32'h00020019;
14'd4758:data <=32'hFFF10019;14'd4759:data <=32'hFFE50020;14'd4760:data <=32'hFFDF002B;
14'd4761:data <=32'hFFDF0035;14'd4762:data <=32'hFFE2003C;14'd4763:data <=32'hFFE60042;
14'd4764:data <=32'hFFEB0046;14'd4765:data <=32'hFFEF004B;14'd4766:data <=32'hFFF40051;
14'd4767:data <=32'hFFFB0056;14'd4768:data <=32'h00050059;14'd4769:data <=32'h0010005A;
14'd4770:data <=32'h001A0058;14'd4771:data <=32'h00220053;14'd4772:data <=32'h0028004D;
14'd4773:data <=32'h002B0049;14'd4774:data <=32'h002D0046;14'd4775:data <=32'h00300046;
14'd4776:data <=32'h00370047;14'd4777:data <=32'h003F0046;14'd4778:data <=32'h004B0043;
14'd4779:data <=32'h0056003B;14'd4780:data <=32'h005D002F;14'd4781:data <=32'h005F001F;
14'd4782:data <=32'h005B0011;14'd4783:data <=32'h00540008;14'd4784:data <=32'h00490004;
14'd4785:data <=32'h00400008;14'd4786:data <=32'h003A0013;14'd4787:data <=32'h003D0020;
14'd4788:data <=32'h0049002C;14'd4789:data <=32'h005D0033;14'd4790:data <=32'h00740034;
14'd4791:data <=32'h008F002C;14'd4792:data <=32'h00A8001D;14'd4793:data <=32'h00C00005;
14'd4794:data <=32'h00D4FFE6;14'd4795:data <=32'h00E4FFBF;14'd4796:data <=32'h00ECFF90;
14'd4797:data <=32'h00E9FF5A;14'd4798:data <=32'h00D7FF21;14'd4799:data <=32'h00B4FEEA;
14'd4800:data <=32'h0033FF56;14'd4801:data <=32'h0026FF35;14'd4802:data <=32'h0024FF1F;
14'd4803:data <=32'h0057FEE1;14'd4804:data <=32'hFFE7FEAA;14'd4805:data <=32'hFFA7FEBB;
14'd4806:data <=32'hFF70FEDB;14'd4807:data <=32'hFF44FF05;14'd4808:data <=32'hFF25FF30;
14'd4809:data <=32'hFF10FF60;14'd4810:data <=32'hFF05FF8D;14'd4811:data <=32'hFF01FFBC;
14'd4812:data <=32'hFF08FFE8;14'd4813:data <=32'hFF170011;14'd4814:data <=32'hFF2E0033;
14'd4815:data <=32'hFF4A004D;14'd4816:data <=32'hFF69005A;14'd4817:data <=32'hFF840060;
14'd4818:data <=32'hFF9B0060;14'd4819:data <=32'hFFAB005D;14'd4820:data <=32'hFFB70059;
14'd4821:data <=32'hFFC00058;14'd4822:data <=32'hFFCA005A;14'd4823:data <=32'hFFD7005C;
14'd4824:data <=32'hFFE6005B;14'd4825:data <=32'hFFF60054;14'd4826:data <=32'h00040048;
14'd4827:data <=32'h000C0037;14'd4828:data <=32'h000D0025;14'd4829:data <=32'h00060015;
14'd4830:data <=32'hFFFA0008;14'd4831:data <=32'hFFEB0004;14'd4832:data <=32'hFFDA0004;
14'd4833:data <=32'hFFCC000C;14'd4834:data <=32'hFFC10017;14'd4835:data <=32'hFFB90025;
14'd4836:data <=32'hFFB30037;14'd4837:data <=32'hFFB20049;14'd4838:data <=32'hFFB6005E;
14'd4839:data <=32'hFFC10073;14'd4840:data <=32'hFFD20086;14'd4841:data <=32'hFFEB0096;
14'd4842:data <=32'h0009009D;14'd4843:data <=32'h0028009C;14'd4844:data <=32'h00450090;
14'd4845:data <=32'h005C007B;14'd4846:data <=32'h006A0061;14'd4847:data <=32'h006C0047;
14'd4848:data <=32'h00650030;14'd4849:data <=32'h00570022;14'd4850:data <=32'h0048001D;
14'd4851:data <=32'h003C0021;14'd4852:data <=32'h0036002C;14'd4853:data <=32'h00370038;
14'd4854:data <=32'h00410045;14'd4855:data <=32'h004F004E;14'd4856:data <=32'h00620052;
14'd4857:data <=32'h00790053;14'd4858:data <=32'h0093004D;14'd4859:data <=32'h00AE003F;
14'd4860:data <=32'h00C90029;14'd4861:data <=32'h00E20009;14'd4862:data <=32'h00F6FFDF;
14'd4863:data <=32'h00FCFFAC;14'd4864:data <=32'h00F6FFEE;14'd4865:data <=32'h0113FFAC;
14'd4866:data <=32'h010DFF7B;14'd4867:data <=32'h00BCFF8B;14'd4868:data <=32'h0073FF43;
14'd4869:data <=32'h0053FF3F;14'd4870:data <=32'h0038FF40;14'd4871:data <=32'h0021FF46;
14'd4872:data <=32'h0011FF4A;14'd4873:data <=32'h0003FF4B;14'd4874:data <=32'hFFF4FF4B;
14'd4875:data <=32'hFFE1FF4C;14'd4876:data <=32'hFFCEFF4C;14'd4877:data <=32'hFFB7FF53;
14'd4878:data <=32'hFFA3FF5D;14'd4879:data <=32'hFF90FF69;14'd4880:data <=32'hFF7FFF77;
14'd4881:data <=32'hFF6EFF88;14'd4882:data <=32'hFF5FFF99;14'd4883:data <=32'hFF4EFFAF;
14'd4884:data <=32'hFF41FFCC;14'd4885:data <=32'hFF38FFEE;14'd4886:data <=32'hFF3B0015;
14'd4887:data <=32'hFF47003B;14'd4888:data <=32'hFF62005E;14'd4889:data <=32'hFF840076;
14'd4890:data <=32'hFFAD0081;14'd4891:data <=32'hFFD4007D;14'd4892:data <=32'hFFF6006E;
14'd4893:data <=32'h00100057;14'd4894:data <=32'h001D003A;14'd4895:data <=32'h0020001D;
14'd4896:data <=32'h001B0004;14'd4897:data <=32'h000FFFEE;14'd4898:data <=32'hFFFCFFDF;
14'd4899:data <=32'hFFE6FFD5;14'd4900:data <=32'hFFCEFFD2;14'd4901:data <=32'hFFB5FFD6;
14'd4902:data <=32'hFF9DFFE2;14'd4903:data <=32'hFF89FFF7;14'd4904:data <=32'hFF7A0013;
14'd4905:data <=32'hFF760033;14'd4906:data <=32'hFF7B0052;14'd4907:data <=32'hFF8A006F;
14'd4908:data <=32'hFF9F0085;14'd4909:data <=32'hFFB70092;14'd4910:data <=32'hFFD00098;
14'd4911:data <=32'hFFE40099;14'd4912:data <=32'hFFF30096;14'd4913:data <=32'h00000094;
14'd4914:data <=32'h00090097;14'd4915:data <=32'h0015009A;14'd4916:data <=32'h002500A0;
14'd4917:data <=32'h003900A4;14'd4918:data <=32'h005000A3;14'd4919:data <=32'h006A009E;
14'd4920:data <=32'h00820091;14'd4921:data <=32'h00980081;14'd4922:data <=32'h00AB006D;
14'd4923:data <=32'h00B90055;14'd4924:data <=32'h00C6003E;14'd4925:data <=32'h00D00023;
14'd4926:data <=32'h00D60004;14'd4927:data <=32'h00D6FFE3;14'd4928:data <=32'h00A100B9;
14'd4929:data <=32'h00EC009E;14'd4930:data <=32'h0117005E;14'd4931:data <=32'h00ACFFBC;
14'd4932:data <=32'h0063FF80;14'd4933:data <=32'h0045FF8A;14'd4934:data <=32'h0031FF9D;
14'd4935:data <=32'h0028FFB2;14'd4936:data <=32'h002DFFC5;14'd4937:data <=32'h003AFFCD;
14'd4938:data <=32'h004AFFCC;14'd4939:data <=32'h0057FFC2;14'd4940:data <=32'h0060FFB0;
14'd4941:data <=32'h0062FF9B;14'd4942:data <=32'h005CFF85;14'd4943:data <=32'h0051FF6F;
14'd4944:data <=32'h0041FF58;14'd4945:data <=32'h0028FF44;14'd4946:data <=32'h0009FF35;
14'd4947:data <=32'hFFE3FF2D;14'd4948:data <=32'hFFB8FF2F;14'd4949:data <=32'hFF8EFF3F;
14'd4950:data <=32'hFF67FF5B;14'd4951:data <=32'hFF4CFF84;14'd4952:data <=32'hFF3FFFB1;
14'd4953:data <=32'hFF40FFDF;14'd4954:data <=32'hFF4E0008;14'd4955:data <=32'hFF690028;
14'd4956:data <=32'hFF85003C;14'd4957:data <=32'hFFA40046;14'd4958:data <=32'hFFBF0046;
14'd4959:data <=32'hFFD60041;14'd4960:data <=32'hFFEA0037;14'd4961:data <=32'hFFF8002A;
14'd4962:data <=32'h0003001B;14'd4963:data <=32'h0009000B;14'd4964:data <=32'h000BFFF7;
14'd4965:data <=32'h0006FFE4;14'd4966:data <=32'hFFFBFFD3;14'd4967:data <=32'hFFEAFFC5;
14'd4968:data <=32'hFFD5FFBE;14'd4969:data <=32'hFFBFFFBE;14'd4970:data <=32'hFFAAFFC3;
14'd4971:data <=32'hFF96FFCD;14'd4972:data <=32'hFF86FFD9;14'd4973:data <=32'hFF78FFE7;
14'd4974:data <=32'hFF6AFFF8;14'd4975:data <=32'hFF5C000B;14'd4976:data <=32'hFF4F0023;
14'd4977:data <=32'hFF440040;14'd4978:data <=32'hFF3D0067;14'd4979:data <=32'hFF410092;
14'd4980:data <=32'hFF5100C1;14'd4981:data <=32'hFF7000ED;14'd4982:data <=32'hFF9C0111;
14'd4983:data <=32'hFFD1012A;14'd4984:data <=32'h000D0133;14'd4985:data <=32'h0047012E;
14'd4986:data <=32'h007E011B;14'd4987:data <=32'h00AF00FD;14'd4988:data <=32'h00D600D7;
14'd4989:data <=32'h00F600A9;14'd4990:data <=32'h010C0077;14'd4991:data <=32'h01140041;
14'd4992:data <=32'h003100AE;14'd4993:data <=32'h006700BB;14'd4994:data <=32'h00AD00AD;
14'd4995:data <=32'h01080015;14'd4996:data <=32'h00C0FFBA;14'd4997:data <=32'h0099FFAC;
14'd4998:data <=32'h0076FFAC;14'd4999:data <=32'h005BFFB6;14'd5000:data <=32'h004DFFC6;
14'd5001:data <=32'h004AFFD4;14'd5002:data <=32'h004DFFDD;14'd5003:data <=32'h0055FFDF;
14'd5004:data <=32'h005DFFDB;14'd5005:data <=32'h0062FFD4;14'd5006:data <=32'h0067FFCA;
14'd5007:data <=32'h0068FFBE;14'd5008:data <=32'h0067FFAF;14'd5009:data <=32'h0064FF9F;
14'd5010:data <=32'h005CFF8C;14'd5011:data <=32'h004EFF79;14'd5012:data <=32'h0038FF69;
14'd5013:data <=32'h001EFF60;14'd5014:data <=32'h0000FF5E;14'd5015:data <=32'hFFE4FF67;
14'd5016:data <=32'hFFCCFF77;14'd5017:data <=32'hFFBDFF8A;14'd5018:data <=32'hFFB5FF9F;
14'd5019:data <=32'hFFB5FFB1;14'd5020:data <=32'hFFB7FFBE;14'd5021:data <=32'hFFB9FFC7;
14'd5022:data <=32'hFFBAFFCD;14'd5023:data <=32'hFFBAFFD3;14'd5024:data <=32'hFFB8FFDB;
14'd5025:data <=32'hFFB7FFE5;14'd5026:data <=32'hFFBBFFF2;14'd5027:data <=32'hFFC2FFFC;
14'd5028:data <=32'hFFCC0004;14'd5029:data <=32'hFFDA0007;14'd5030:data <=32'hFFE80005;
14'd5031:data <=32'hFFF3FFFF;14'd5032:data <=32'hFFFCFFF4;14'd5033:data <=32'h0002FFE6;
14'd5034:data <=32'h0003FFD6;14'd5035:data <=32'h0000FFC6;14'd5036:data <=32'hFFFAFFB4;
14'd5037:data <=32'hFFEBFFA0;14'd5038:data <=32'hFFD6FF8F;14'd5039:data <=32'hFFB8FF80;
14'd5040:data <=32'hFF91FF79;14'd5041:data <=32'hFF64FF7F;14'd5042:data <=32'hFF35FF93;
14'd5043:data <=32'hFF0AFFB9;14'd5044:data <=32'hFEE9FFEC;14'd5045:data <=32'hFEDA002B;
14'd5046:data <=32'hFEDB006D;14'd5047:data <=32'hFEEF00AD;14'd5048:data <=32'hFF1400E6;
14'd5049:data <=32'hFF430113;14'd5050:data <=32'hFF7B0132;14'd5051:data <=32'hFFB60144;
14'd5052:data <=32'hFFF40149;14'd5053:data <=32'h002F0141;14'd5054:data <=32'h0068012D;
14'd5055:data <=32'h0099010E;14'd5056:data <=32'h003300D2;14'd5057:data <=32'h005C00D9;
14'd5058:data <=32'h008500E4;14'd5059:data <=32'h00AF00FB;14'd5060:data <=32'h009A00A0;
14'd5061:data <=32'h009F0086;14'd5062:data <=32'h00A30074;14'd5063:data <=32'h00A60063;
14'd5064:data <=32'h00AC0056;14'd5065:data <=32'h00B70045;14'd5066:data <=32'h00C2002F;
14'd5067:data <=32'h00C80015;14'd5068:data <=32'h00C9FFF7;14'd5069:data <=32'h00C1FFD7;
14'd5070:data <=32'h00B1FFBA;14'd5071:data <=32'h009DFFA5;14'd5072:data <=32'h0086FF95;
14'd5073:data <=32'h006FFF8C;14'd5074:data <=32'h0058FF86;14'd5075:data <=32'h0042FF85;
14'd5076:data <=32'h002CFF86;14'd5077:data <=32'h0017FF8C;14'd5078:data <=32'h0004FF98;
14'd5079:data <=32'hFFF7FFA9;14'd5080:data <=32'hFFF0FFBC;14'd5081:data <=32'hFFF2FFCF;
14'd5082:data <=32'hFFFBFFDF;14'd5083:data <=32'h000AFFE7;14'd5084:data <=32'h001BFFE6;
14'd5085:data <=32'h0028FFDC;14'd5086:data <=32'h002FFFCC;14'd5087:data <=32'h002DFFBA;
14'd5088:data <=32'h0023FFAB;14'd5089:data <=32'h0014FFA1;14'd5090:data <=32'h0001FF9E;
14'd5091:data <=32'hFFF2FFA2;14'd5092:data <=32'hFFE4FFA9;14'd5093:data <=32'hFFDDFFB4;
14'd5094:data <=32'hFFD9FFC0;14'd5095:data <=32'hFFD9FFC9;14'd5096:data <=32'hFFDCFFD2;
14'd5097:data <=32'hFFE1FFD7;14'd5098:data <=32'hFFE8FFD9;14'd5099:data <=32'hFFF1FFD9;
14'd5100:data <=32'hFFFAFFD2;14'd5101:data <=32'h0002FFC7;14'd5102:data <=32'h0005FFB5;
14'd5103:data <=32'h0001FF9F;14'd5104:data <=32'hFFF2FF88;14'd5105:data <=32'hFFDAFF73;
14'd5106:data <=32'hFFB7FF67;14'd5107:data <=32'hFF8FFF66;14'd5108:data <=32'hFF65FF75;
14'd5109:data <=32'hFF40FF8E;14'd5110:data <=32'hFF25FFB2;14'd5111:data <=32'hFF14FFDA;
14'd5112:data <=32'hFF0E0004;14'd5113:data <=32'hFF11002C;14'd5114:data <=32'hFF1A0050;
14'd5115:data <=32'hFF280070;14'd5116:data <=32'hFF39008E;14'd5117:data <=32'hFF4F00A8;
14'd5118:data <=32'hFF6800C0;14'd5119:data <=32'hFF8600D5;14'd5120:data <=32'hFF93011A;
14'd5121:data <=32'hFFC60136;14'd5122:data <=32'hFFEA0137;14'd5123:data <=32'hFF9700F1;
14'd5124:data <=32'hFF8900C8;14'd5125:data <=32'hFF9D00E1;14'd5126:data <=32'hFFB900F9;
14'd5127:data <=32'hFFDD010F;14'd5128:data <=32'h000A0120;14'd5129:data <=32'h00410126;
14'd5130:data <=32'h007C011C;14'd5131:data <=32'h00B40101;14'd5132:data <=32'h00E400D6;
14'd5133:data <=32'h010600A1;14'd5134:data <=32'h01170064;14'd5135:data <=32'h01170028;
14'd5136:data <=32'h010BFFF2;14'd5137:data <=32'h00F3FFC3;14'd5138:data <=32'h00D3FF9D;
14'd5139:data <=32'h00AEFF81;14'd5140:data <=32'h0085FF6E;14'd5141:data <=32'h005AFF67;
14'd5142:data <=32'h002FFF6B;14'd5143:data <=32'h0008FF7C;14'd5144:data <=32'hFFEAFF96;
14'd5145:data <=32'hFFD8FFB8;14'd5146:data <=32'hFFD4FFDB;14'd5147:data <=32'hFFDEFFFB;
14'd5148:data <=32'hFFF20012;14'd5149:data <=32'h000A001E;14'd5150:data <=32'h0022001F;
14'd5151:data <=32'h00380017;14'd5152:data <=32'h00460009;14'd5153:data <=32'h004EFFF9;
14'd5154:data <=32'h0051FFEB;14'd5155:data <=32'h0051FFDF;14'd5156:data <=32'h004FFFD4;
14'd5157:data <=32'h004DFFC9;14'd5158:data <=32'h004BFFBF;14'd5159:data <=32'h0048FFB3;
14'd5160:data <=32'h0042FFA8;14'd5161:data <=32'h0039FF9E;14'd5162:data <=32'h002FFF95;
14'd5163:data <=32'h0024FF8E;14'd5164:data <=32'h0019FF89;14'd5165:data <=32'h000EFF83;
14'd5166:data <=32'h0004FF7F;14'd5167:data <=32'hFFF8FF7A;14'd5168:data <=32'hFFEAFF75;
14'd5169:data <=32'hFFD8FF70;14'd5170:data <=32'hFFC2FF6F;14'd5171:data <=32'hFFA9FF74;
14'd5172:data <=32'hFF92FF82;14'd5173:data <=32'hFF80FF94;14'd5174:data <=32'hFF74FFAD;
14'd5175:data <=32'hFF71FFC5;14'd5176:data <=32'hFF75FFD9;14'd5177:data <=32'hFF7EFFE7;
14'd5178:data <=32'hFF86FFEE;14'd5179:data <=32'hFF8BFFEE;14'd5180:data <=32'hFF8BFFEB;
14'd5181:data <=32'hFF83FFEB;14'd5182:data <=32'hFF78FFED;14'd5183:data <=32'hFF69FFF5;
14'd5184:data <=32'hFEF1005E;14'd5185:data <=32'hFEFA0094;14'd5186:data <=32'hFF2000AD;
14'd5187:data <=32'hFF5A0021;14'd5188:data <=32'hFF27FFFD;14'd5189:data <=32'hFF120024;
14'd5190:data <=32'hFF060053;14'd5191:data <=32'hFF08008A;14'd5192:data <=32'hFF1A00C3;
14'd5193:data <=32'hFF3E00FA;14'd5194:data <=32'hFF730125;14'd5195:data <=32'hFFB5013F;
14'd5196:data <=32'hFFF90145;14'd5197:data <=32'h003B0139;14'd5198:data <=32'h0074011C;
14'd5199:data <=32'h00A100F5;14'd5200:data <=32'h00C200C9;14'd5201:data <=32'h00D70099;
14'd5202:data <=32'h00E10068;14'd5203:data <=32'h00E2003A;14'd5204:data <=32'h00D8000E;
14'd5205:data <=32'h00C5FFE7;14'd5206:data <=32'h00A9FFC5;14'd5207:data <=32'h0087FFAF;
14'd5208:data <=32'h0063FFA4;14'd5209:data <=32'h0040FFA5;14'd5210:data <=32'h0024FFB1;
14'd5211:data <=32'h000FFFC2;14'd5212:data <=32'h0004FFD5;14'd5213:data <=32'hFFFFFFE7;
14'd5214:data <=32'hFFFFFFF4;14'd5215:data <=32'h0002FFFF;14'd5216:data <=32'h00040009;
14'd5217:data <=32'h00070012;14'd5218:data <=32'h000B001E;14'd5219:data <=32'h0013002A;
14'd5220:data <=32'h00210036;14'd5221:data <=32'h0035003E;14'd5222:data <=32'h004E0040;
14'd5223:data <=32'h0068003B;14'd5224:data <=32'h0082002B;14'd5225:data <=32'h00980014;
14'd5226:data <=32'h00A8FFF7;14'd5227:data <=32'h00AEFFD5;14'd5228:data <=32'h00AEFFB3;
14'd5229:data <=32'h00A5FF90;14'd5230:data <=32'h0096FF6F;14'd5231:data <=32'h0080FF51;
14'd5232:data <=32'h0062FF38;14'd5233:data <=32'h003EFF23;14'd5234:data <=32'h0014FF18;
14'd5235:data <=32'hFFE7FF18;14'd5236:data <=32'hFFBBFF25;14'd5237:data <=32'hFF95FF3E;
14'd5238:data <=32'hFF79FF62;14'd5239:data <=32'hFF6DFF89;14'd5240:data <=32'hFF6DFFAF;
14'd5241:data <=32'hFF79FFCD;14'd5242:data <=32'hFF8DFFE0;14'd5243:data <=32'hFFA2FFE7;
14'd5244:data <=32'hFFB2FFE4;14'd5245:data <=32'hFFBCFFDA;14'd5246:data <=32'hFFBEFFCD;
14'd5247:data <=32'hFFB9FFC0;14'd5248:data <=32'hFF70FF9C;14'd5249:data <=32'hFF53FFA7;
14'd5250:data <=32'hFF4CFFC8;14'd5251:data <=32'hFF93FFED;14'd5252:data <=32'hFF65FFB3;
14'd5253:data <=32'hFF4DFFC2;14'd5254:data <=32'hFF38FFDA;14'd5255:data <=32'hFF26FFF8;
14'd5256:data <=32'hFF1C0021;14'd5257:data <=32'hFF1F004D;14'd5258:data <=32'hFF2F0078;
14'd5259:data <=32'hFF4B009C;14'd5260:data <=32'hFF6F00B5;14'd5261:data <=32'hFF9500C3;
14'd5262:data <=32'hFFB800C7;14'd5263:data <=32'hFFD800C3;14'd5264:data <=32'hFFF100BC;
14'd5265:data <=32'h000600B4;14'd5266:data <=32'h001900AA;14'd5267:data <=32'h002C00A1;
14'd5268:data <=32'h003F0094;14'd5269:data <=32'h004E0085;14'd5270:data <=32'h005C0072;
14'd5271:data <=32'h0064005F;14'd5272:data <=32'h0066004D;14'd5273:data <=32'h0066003B;
14'd5274:data <=32'h0064002D;14'd5275:data <=32'h00610020;14'd5276:data <=32'h005F0014;
14'd5277:data <=32'h005C0006;14'd5278:data <=32'h0055FFF8;14'd5279:data <=32'h0049FFE9;
14'd5280:data <=32'h0036FFDE;14'd5281:data <=32'h0021FFD9;14'd5282:data <=32'h0007FFDE;
14'd5283:data <=32'hFFF0FFEC;14'd5284:data <=32'hFFE10005;14'd5285:data <=32'hFFDB0023;
14'd5286:data <=32'hFFE20044;14'd5287:data <=32'hFFF60060;14'd5288:data <=32'h00120075;
14'd5289:data <=32'h00350080;14'd5290:data <=32'h005B007F;14'd5291:data <=32'h007F0076;
14'd5292:data <=32'h00A10062;14'd5293:data <=32'h00BE0045;14'd5294:data <=32'h00D50023;
14'd5295:data <=32'h00E2FFFB;14'd5296:data <=32'h00E7FFCE;14'd5297:data <=32'h00E0FF9F;
14'd5298:data <=32'h00CEFF72;14'd5299:data <=32'h00AFFF4D;14'd5300:data <=32'h0088FF30;
14'd5301:data <=32'h005CFF22;14'd5302:data <=32'h0031FF1F;14'd5303:data <=32'h000CFF28;
14'd5304:data <=32'hFFEFFF39;14'd5305:data <=32'hFFDCFF4B;14'd5306:data <=32'hFFD1FF5B;
14'd5307:data <=32'hFFCAFF66;14'd5308:data <=32'hFFC5FF6B;14'd5309:data <=32'hFFBDFF6E;
14'd5310:data <=32'hFFB0FF71;14'd5311:data <=32'hFFA2FF75;14'd5312:data <=32'hFFECFFC7;
14'd5313:data <=32'hFFEEFFAE;14'd5314:data <=32'hFFD8FF9E;14'd5315:data <=32'hFF65FF9F;
14'd5316:data <=32'hFF3BFF7A;14'd5317:data <=32'hFF2AFF9A;14'd5318:data <=32'hFF1FFFBD;
14'd5319:data <=32'hFF1BFFE2;14'd5320:data <=32'hFF1E0009;14'd5321:data <=32'hFF2B002F;
14'd5322:data <=32'hFF430051;14'd5323:data <=32'hFF62006A;14'd5324:data <=32'hFF850076;
14'd5325:data <=32'hFFA80075;14'd5326:data <=32'hFFC3006A;14'd5327:data <=32'hFFD50058;
14'd5328:data <=32'hFFDB0046;14'd5329:data <=32'hFFD8003A;14'd5330:data <=32'hFFD10033;
14'd5331:data <=32'hFFC70032;14'd5332:data <=32'hFFBF003A;14'd5333:data <=32'hFFBE0044;
14'd5334:data <=32'hFFC00050;14'd5335:data <=32'hFFC5005C;14'd5336:data <=32'hFFCC0068;
14'd5337:data <=32'hFFD80073;14'd5338:data <=32'hFFE7007B;14'd5339:data <=32'hFFFA0084;
14'd5340:data <=32'h00120085;14'd5341:data <=32'h002B007F;14'd5342:data <=32'h00410070;
14'd5343:data <=32'h00530059;14'd5344:data <=32'h005A003E;14'd5345:data <=32'h00570021;
14'd5346:data <=32'h0049000A;14'd5347:data <=32'h0033FFFA;14'd5348:data <=32'h001CFFF6;
14'd5349:data <=32'h0004FFFB;14'd5350:data <=32'hFFF4000A;14'd5351:data <=32'hFFE9001D;
14'd5352:data <=32'hFFE80034;14'd5353:data <=32'hFFED0047;14'd5354:data <=32'hFFFA0059;
14'd5355:data <=32'h00090067;14'd5356:data <=32'h001B0071;14'd5357:data <=32'h00300077;
14'd5358:data <=32'h0048007B;14'd5359:data <=32'h00610078;14'd5360:data <=32'h007C006F;
14'd5361:data <=32'h00940061;14'd5362:data <=32'h00AA004B;14'd5363:data <=32'h00BA0031;
14'd5364:data <=32'h00C30015;14'd5365:data <=32'h00C7FFFB;14'd5366:data <=32'h00C7FFE1;
14'd5367:data <=32'h00C5FFCB;14'd5368:data <=32'h00C4FFB6;14'd5369:data <=32'h00C3FF9E;
14'd5370:data <=32'h00C2FF82;14'd5371:data <=32'h00BCFF60;14'd5372:data <=32'h00ADFF3A;
14'd5373:data <=32'h0094FF15;14'd5374:data <=32'h006EFEF3;14'd5375:data <=32'h003EFEDB;
14'd5376:data <=32'hFFEAFFBB;14'd5377:data <=32'hFFFAFFB3;14'd5378:data <=32'h000AFF91;
14'd5379:data <=32'hFFE5FEE7;14'd5380:data <=32'hFF93FEB8;14'd5381:data <=32'hFF5AFED8;
14'd5382:data <=32'hFF2BFF04;14'd5383:data <=32'hFF07FF39;14'd5384:data <=32'hFEEFFF74;
14'd5385:data <=32'hFEE8FFB4;14'd5386:data <=32'hFEF2FFF0;14'd5387:data <=32'hFF0D0026;
14'd5388:data <=32'hFF35004F;14'd5389:data <=32'hFF630066;14'd5390:data <=32'hFF91006B;
14'd5391:data <=32'hFFB80061;14'd5392:data <=32'hFFD2004F;14'd5393:data <=32'hFFE1003A;
14'd5394:data <=32'hFFE50025;14'd5395:data <=32'hFFE20014;14'd5396:data <=32'hFFDA000B;
14'd5397:data <=32'hFFD10005;14'd5398:data <=32'hFFC70004;14'd5399:data <=32'hFFBD0006;
14'd5400:data <=32'hFFB4000C;14'd5401:data <=32'hFFAC0016;14'd5402:data <=32'hFFA60022;
14'd5403:data <=32'hFFA60033;14'd5404:data <=32'hFFAA0044;14'd5405:data <=32'hFFB50054;
14'd5406:data <=32'hFFC6005E;14'd5407:data <=32'hFFD80063;14'd5408:data <=32'hFFE90060;
14'd5409:data <=32'hFFF60059;14'd5410:data <=32'hFFFD0050;14'd5411:data <=32'hFFFF0048;
14'd5412:data <=32'hFFFD0043;14'd5413:data <=32'hFFF90043;14'd5414:data <=32'hFFFA0046;
14'd5415:data <=32'hFFFD004A;14'd5416:data <=32'h0003004E;14'd5417:data <=32'h000A004F;
14'd5418:data <=32'h0012004C;14'd5419:data <=32'h00180046;14'd5420:data <=32'h00190040;
14'd5421:data <=32'h0016003B;14'd5422:data <=32'h0011003B;14'd5423:data <=32'h000C0040;
14'd5424:data <=32'h000A0047;14'd5425:data <=32'h000C0051;14'd5426:data <=32'h0010005E;
14'd5427:data <=32'h0018006A;14'd5428:data <=32'h00260076;14'd5429:data <=32'h00340082;
14'd5430:data <=32'h004B008C;14'd5431:data <=32'h00670096;14'd5432:data <=32'h008B0099;
14'd5433:data <=32'h00B50093;14'd5434:data <=32'h00E40080;14'd5435:data <=32'h0111005C;
14'd5436:data <=32'h01360028;14'd5437:data <=32'h014DFFE6;14'd5438:data <=32'h014FFF9E;
14'd5439:data <=32'h013EFF55;14'd5440:data <=32'h0079FF99;14'd5441:data <=32'h0082FF82;
14'd5442:data <=32'h0097FF73;14'd5443:data <=32'h00F0FF38;14'd5444:data <=32'h00A9FED3;
14'd5445:data <=32'h006CFEBF;14'd5446:data <=32'h002EFEB8;14'd5447:data <=32'hFFF2FEBF;
14'd5448:data <=32'hFFB9FED3;14'd5449:data <=32'hFF87FEF5;14'd5450:data <=32'hFF61FF20;
14'd5451:data <=32'hFF4BFF50;14'd5452:data <=32'hFF43FF80;14'd5453:data <=32'hFF48FFA9;
14'd5454:data <=32'hFF57FFC8;14'd5455:data <=32'hFF67FFDF;14'd5456:data <=32'hFF76FFEC;
14'd5457:data <=32'hFF81FFF5;14'd5458:data <=32'hFF88FFFD;14'd5459:data <=32'hFF8F0006;
14'd5460:data <=32'hFF950010;14'd5461:data <=32'hFF9F001A;14'd5462:data <=32'hFFAA0021;
14'd5463:data <=32'hFFBA0025;14'd5464:data <=32'hFFC60024;14'd5465:data <=32'hFFCF001F;
14'd5466:data <=32'hFFD50019;14'd5467:data <=32'hFFD70013;14'd5468:data <=32'hFFD9000E;
14'd5469:data <=32'hFFD8000A;14'd5470:data <=32'hFFD80006;14'd5471:data <=32'hFFD60002;
14'd5472:data <=32'hFFD1FFFD;14'd5473:data <=32'hFFC9FFF8;14'd5474:data <=32'hFFBDFFF7;
14'd5475:data <=32'hFFAEFFFC;14'd5476:data <=32'hFF9E0006;14'd5477:data <=32'hFF930019;
14'd5478:data <=32'hFF8E0031;14'd5479:data <=32'hFF91004B;14'd5480:data <=32'hFF9F0063;
14'd5481:data <=32'hFFB50075;14'd5482:data <=32'hFFCE007F;14'd5483:data <=32'hFFE8007F;
14'd5484:data <=32'hFFFC0077;14'd5485:data <=32'h000B0069;14'd5486:data <=32'h0012005B;
14'd5487:data <=32'h0013004E;14'd5488:data <=32'h000F0044;14'd5489:data <=32'h0008003F;
14'd5490:data <=32'hFFFF003E;14'd5491:data <=32'hFFF70042;14'd5492:data <=32'hFFEF004A;
14'd5493:data <=32'hFFE9005A;14'd5494:data <=32'hFFE7006E;14'd5495:data <=32'hFFED0088;
14'd5496:data <=32'hFFFD00A3;14'd5497:data <=32'h001A00BD;14'd5498:data <=32'h004300CF;
14'd5499:data <=32'h007500D6;14'd5500:data <=32'h00AC00CA;14'd5501:data <=32'h00DF00AE;
14'd5502:data <=32'h01090082;14'd5503:data <=32'h0125004C;14'd5504:data <=32'h00E80069;
14'd5505:data <=32'h01170044;14'd5506:data <=32'h012A0025;14'd5507:data <=32'h00F70025;
14'd5508:data <=32'h00DFFFC2;14'd5509:data <=32'h00D2FFA7;14'd5510:data <=32'h00C2FF8D;
14'd5511:data <=32'h00AFFF78;14'd5512:data <=32'h0099FF64;14'd5513:data <=32'h007FFF56;
14'd5514:data <=32'h0066FF4D;14'd5515:data <=32'h004EFF49;14'd5516:data <=32'h003AFF47;
14'd5517:data <=32'h0029FF46;14'd5518:data <=32'h0017FF43;14'd5519:data <=32'h0004FF3D;
14'd5520:data <=32'hFFECFF39;14'd5521:data <=32'hFFCDFF38;14'd5522:data <=32'hFFAAFF40;
14'd5523:data <=32'hFF88FF51;14'd5524:data <=32'hFF6BFF6E;14'd5525:data <=32'hFF57FF93;
14'd5526:data <=32'hFF50FFBC;14'd5527:data <=32'hFF55FFE4;14'd5528:data <=32'hFF640005;
14'd5529:data <=32'hFF780020;14'd5530:data <=32'hFF920032;14'd5531:data <=32'hFFAE003B;
14'd5532:data <=32'hFFC8003E;14'd5533:data <=32'hFFE2003A;14'd5534:data <=32'hFFF8002E;
14'd5535:data <=32'h000B001C;14'd5536:data <=32'h00170004;14'd5537:data <=32'h0019FFE9;
14'd5538:data <=32'h0011FFCE;14'd5539:data <=32'hFFFDFFB6;14'd5540:data <=32'hFFE1FFA8;
14'd5541:data <=32'hFFC1FFA5;14'd5542:data <=32'hFFA2FFAC;14'd5543:data <=32'hFF87FFBF;
14'd5544:data <=32'hFF76FFD9;14'd5545:data <=32'hFF6DFFF5;14'd5546:data <=32'hFF6E0010;
14'd5547:data <=32'hFF750027;14'd5548:data <=32'hFF7E0038;14'd5549:data <=32'hFF890045;
14'd5550:data <=32'hFF92004F;14'd5551:data <=32'hFF990056;14'd5552:data <=32'hFFA0005F;
14'd5553:data <=32'hFFA8006A;14'd5554:data <=32'hFFB00073;14'd5555:data <=32'hFFBA007C;
14'd5556:data <=32'hFFC30083;14'd5557:data <=32'hFFCE008B;14'd5558:data <=32'hFFD80093;
14'd5559:data <=32'hFFE2009D;14'd5560:data <=32'hFFF000A8;14'd5561:data <=32'h000300B5;
14'd5562:data <=32'h001D00BE;14'd5563:data <=32'h003D00C3;14'd5564:data <=32'h006000BE;
14'd5565:data <=32'h008200AD;14'd5566:data <=32'h009E0096;14'd5567:data <=32'h00B00075;
14'd5568:data <=32'h0037010C;14'd5569:data <=32'h0081011A;14'd5570:data <=32'h00BC00FC;
14'd5571:data <=32'h00910054;14'd5572:data <=32'h00770009;14'd5573:data <=32'h006B000A;
14'd5574:data <=32'h0066000E;14'd5575:data <=32'h00680014;14'd5576:data <=32'h006E0016;
14'd5577:data <=32'h00760015;14'd5578:data <=32'h00810012;14'd5579:data <=32'h008F000B;
14'd5580:data <=32'h009FFFFF;14'd5581:data <=32'h00B0FFEC;14'd5582:data <=32'h00BDFFCF;
14'd5583:data <=32'h00C2FFA9;14'd5584:data <=32'h00BDFF7F;14'd5585:data <=32'h00A8FF54;
14'd5586:data <=32'h0085FF2E;14'd5587:data <=32'h0056FF15;14'd5588:data <=32'h0022FF0A;
14'd5589:data <=32'hFFEDFF10;14'd5590:data <=32'hFFC0FF25;14'd5591:data <=32'hFF9BFF44;
14'd5592:data <=32'hFF82FF68;14'd5593:data <=32'hFF74FF8E;14'd5594:data <=32'hFF6FFFB2;
14'd5595:data <=32'hFF74FFD4;14'd5596:data <=32'hFF80FFF3;14'd5597:data <=32'hFF92000D;
14'd5598:data <=32'hFFA90020;14'd5599:data <=32'hFFC5002C;14'd5600:data <=32'hFFE2002D;
14'd5601:data <=32'hFFFE0026;14'd5602:data <=32'h00130014;14'd5603:data <=32'h0022FFFD;
14'd5604:data <=32'h0025FFE3;14'd5605:data <=32'h0020FFCB;14'd5606:data <=32'h0014FFB7;
14'd5607:data <=32'h0005FFAA;14'd5608:data <=32'hFFF3FFA1;14'd5609:data <=32'hFFE3FF9D;
14'd5610:data <=32'hFFD3FF99;14'd5611:data <=32'hFFC3FF96;14'd5612:data <=32'hFFB1FF93;
14'd5613:data <=32'hFF9BFF93;14'd5614:data <=32'hFF80FF96;14'd5615:data <=32'hFF63FFA2;
14'd5616:data <=32'hFF45FFB6;14'd5617:data <=32'hFF2CFFD4;14'd5618:data <=32'hFF19FFF9;
14'd5619:data <=32'hFF110023;14'd5620:data <=32'hFF11004F;14'd5621:data <=32'hFF1B007A;
14'd5622:data <=32'hFF2E00A4;14'd5623:data <=32'hFF4900C9;14'd5624:data <=32'hFF6B00E9;
14'd5625:data <=32'hFF940104;14'd5626:data <=32'hFFC40115;14'd5627:data <=32'hFFFA011B;
14'd5628:data <=32'h00310115;14'd5629:data <=32'h006300FE;14'd5630:data <=32'h008E00DA;
14'd5631:data <=32'h00AA00AD;14'd5632:data <=32'hFFAF00B8;14'd5633:data <=32'hFFD100E3;
14'd5634:data <=32'h001000FC;14'd5635:data <=32'h009A008E;14'd5636:data <=32'h00800031;
14'd5637:data <=32'h006D0023;14'd5638:data <=32'h005C001F;14'd5639:data <=32'h00500023;
14'd5640:data <=32'h00480027;14'd5641:data <=32'h0046002F;14'd5642:data <=32'h00480037;
14'd5643:data <=32'h0050003F;14'd5644:data <=32'h005D0045;14'd5645:data <=32'h00710048;
14'd5646:data <=32'h00880041;14'd5647:data <=32'h00A10031;14'd5648:data <=32'h00B50015;
14'd5649:data <=32'h00C0FFF1;14'd5650:data <=32'h00BFFFCA;14'd5651:data <=32'h00B0FFA6;
14'd5652:data <=32'h0098FF88;14'd5653:data <=32'h007AFF74;14'd5654:data <=32'h005AFF6B;
14'd5655:data <=32'h003EFF69;14'd5656:data <=32'h0025FF6D;14'd5657:data <=32'h0010FF73;
14'd5658:data <=32'hFFFFFF7C;14'd5659:data <=32'hFFEFFF86;14'd5660:data <=32'hFFE1FF91;
14'd5661:data <=32'hFFD6FF9E;14'd5662:data <=32'hFFCDFFAF;14'd5663:data <=32'hFFC8FFC0;
14'd5664:data <=32'hFFCAFFD0;14'd5665:data <=32'hFFD0FFE0;14'd5666:data <=32'hFFD9FFEA;
14'd5667:data <=32'hFFE3FFF1;14'd5668:data <=32'hFFEEFFF6;14'd5669:data <=32'hFFF7FFF6;
14'd5670:data <=32'h0001FFF5;14'd5671:data <=32'h000AFFF4;14'd5672:data <=32'h0017FFF0;
14'd5673:data <=32'h0025FFE9;14'd5674:data <=32'h0032FFDA;14'd5675:data <=32'h003EFFC4;
14'd5676:data <=32'h0043FFA6;14'd5677:data <=32'h003DFF83;14'd5678:data <=32'h002AFF5F;
14'd5679:data <=32'h0008FF3F;14'd5680:data <=32'hFFDCFF2A;14'd5681:data <=32'hFFA6FF21;
14'd5682:data <=32'hFF70FF28;14'd5683:data <=32'hFF3BFF3E;14'd5684:data <=32'hFF0DFF62;
14'd5685:data <=32'hFEE9FF90;14'd5686:data <=32'hFECEFFC6;14'd5687:data <=32'hFEC10000;
14'd5688:data <=32'hFEC0003E;14'd5689:data <=32'hFECE007B;14'd5690:data <=32'hFEE900B7;
14'd5691:data <=32'hFF1500EA;14'd5692:data <=32'hFF4B010F;14'd5693:data <=32'hFF8A0125;
14'd5694:data <=32'hFFC90129;14'd5695:data <=32'h00030119;14'd5696:data <=32'hFFB500A5;
14'd5697:data <=32'hFFC600BA;14'd5698:data <=32'hFFD700DC;14'd5699:data <=32'h00020111;
14'd5700:data <=32'h000E00C2;14'd5701:data <=32'h001E00BB;14'd5702:data <=32'h002D00B4;
14'd5703:data <=32'h003E00AF;14'd5704:data <=32'h005000A6;14'd5705:data <=32'h00610098;
14'd5706:data <=32'h006F0089;14'd5707:data <=32'h007A0079;14'd5708:data <=32'h00840068;
14'd5709:data <=32'h008C0059;14'd5710:data <=32'h00950048;14'd5711:data <=32'h009B0035;
14'd5712:data <=32'h00A0001D;14'd5713:data <=32'h009F0003;14'd5714:data <=32'h0096FFEA;
14'd5715:data <=32'h0085FFD3;14'd5716:data <=32'h006FFFC5;14'd5717:data <=32'h0057FFBF;
14'd5718:data <=32'h0042FFC4;14'd5719:data <=32'h0033FFCE;14'd5720:data <=32'h002DFFDB;
14'd5721:data <=32'h002FFFE5;14'd5722:data <=32'h0035FFEA;14'd5723:data <=32'h003DFFEB;
14'd5724:data <=32'h0043FFE5;14'd5725:data <=32'h0046FFDB;14'd5726:data <=32'h0045FFD2;
14'd5727:data <=32'h0041FFC9;14'd5728:data <=32'h0039FFC0;14'd5729:data <=32'h0031FFBB;
14'd5730:data <=32'h0029FFB5;14'd5731:data <=32'h001EFFB3;14'd5732:data <=32'h0013FFB4;
14'd5733:data <=32'h0008FFB7;14'd5734:data <=32'hFFFDFFBF;14'd5735:data <=32'hFFF7FFCD;
14'd5736:data <=32'hFFF7FFDC;14'd5737:data <=32'hFFFFFFEB;14'd5738:data <=32'h0010FFF6;
14'd5739:data <=32'h0025FFF8;14'd5740:data <=32'h003DFFF0;14'd5741:data <=32'h0053FFDB;
14'd5742:data <=32'h0060FFBE;14'd5743:data <=32'h0062FF98;14'd5744:data <=32'h0057FF74;
14'd5745:data <=32'h003FFF53;14'd5746:data <=32'h001DFF39;14'd5747:data <=32'hFFF7FF29;
14'd5748:data <=32'hFFCEFF23;14'd5749:data <=32'hFFA4FF26;14'd5750:data <=32'hFF7BFF32;
14'd5751:data <=32'hFF55FF45;14'd5752:data <=32'hFF32FF60;14'd5753:data <=32'hFF15FF82;
14'd5754:data <=32'hFF00FFAC;14'd5755:data <=32'hFEF4FFDA;14'd5756:data <=32'hFEF40008;
14'd5757:data <=32'hFEFF0033;14'd5758:data <=32'hFF120057;14'd5759:data <=32'hFF2A0072;
14'd5760:data <=32'hFF3800A6;14'd5761:data <=32'hFF5000C5;14'd5762:data <=32'hFF5D00CE;
14'd5763:data <=32'hFF150086;14'd5764:data <=32'hFF110065;14'd5765:data <=32'hFF180091;
14'd5766:data <=32'hFF2A00BE;14'd5767:data <=32'hFF4900E8;14'd5768:data <=32'hFF74010B;
14'd5769:data <=32'hFFA90121;14'd5770:data <=32'hFFE00129;14'd5771:data <=32'h00160125;
14'd5772:data <=32'h00490115;14'd5773:data <=32'h007700FD;14'd5774:data <=32'h009D00DC;
14'd5775:data <=32'h00BD00B4;14'd5776:data <=32'h00D30085;14'd5777:data <=32'h00DC0052;
14'd5778:data <=32'h00D6001E;14'd5779:data <=32'h00C3FFEF;14'd5780:data <=32'h00A3FFCA;
14'd5781:data <=32'h007BFFB4;14'd5782:data <=32'h0050FFAD;14'd5783:data <=32'h002BFFB5;
14'd5784:data <=32'h000FFFC8;14'd5785:data <=32'hFFFFFFE0;14'd5786:data <=32'hFFFBFFF9;
14'd5787:data <=32'hFFFE000F;14'd5788:data <=32'h0009001E;14'd5789:data <=32'h00170028;
14'd5790:data <=32'h0026002D;14'd5791:data <=32'h0032002C;14'd5792:data <=32'h0041002A;
14'd5793:data <=32'h004D0023;14'd5794:data <=32'h00580019;14'd5795:data <=32'h0060000D;
14'd5796:data <=32'h0064FFFF;14'd5797:data <=32'h0065FFEF;14'd5798:data <=32'h0061FFE1;
14'd5799:data <=32'h0058FFD8;14'd5800:data <=32'h004FFFD2;14'd5801:data <=32'h004AFFD1;
14'd5802:data <=32'h0047FFD1;14'd5803:data <=32'h0049FFD2;14'd5804:data <=32'h004FFFCE;
14'd5805:data <=32'h0056FFC5;14'd5806:data <=32'h005AFFB6;14'd5807:data <=32'h0058FFA4;
14'd5808:data <=32'h0050FF8F;14'd5809:data <=32'h0041FF7F;14'd5810:data <=32'h002DFF73;
14'd5811:data <=32'h001AFF6F;14'd5812:data <=32'h0007FF6F;14'd5813:data <=32'hFFF8FF72;
14'd5814:data <=32'hFFEBFF75;14'd5815:data <=32'hFFE2FF78;14'd5816:data <=32'hFFD8FF7A;
14'd5817:data <=32'hFFCEFF7A;14'd5818:data <=32'hFFC2FF7A;14'd5819:data <=32'hFFB6FF7B;
14'd5820:data <=32'hFFA9FF7F;14'd5821:data <=32'hFF9CFF81;14'd5822:data <=32'hFF8EFF83;
14'd5823:data <=32'hFF7FFF84;14'd5824:data <=32'hFEFAFFCF;14'd5825:data <=32'hFEEDFFF4;
14'd5826:data <=32'hFEFE0009;14'd5827:data <=32'hFF4CFF8F;14'd5828:data <=32'hFF1CFF60;
14'd5829:data <=32'hFEEEFF87;14'd5830:data <=32'hFECBFFBD;14'd5831:data <=32'hFEB7FFFF;
14'd5832:data <=32'hFEB70044;14'd5833:data <=32'hFECB0085;14'd5834:data <=32'hFEEC00BE;
14'd5835:data <=32'hFF1A00ED;14'd5836:data <=32'hFF4F010E;14'd5837:data <=32'hFF870124;
14'd5838:data <=32'hFFC3012E;14'd5839:data <=32'hFFFF0129;14'd5840:data <=32'h00380117;
14'd5841:data <=32'h006A00F7;14'd5842:data <=32'h009000CB;14'd5843:data <=32'h00A9009A;
14'd5844:data <=32'h00AF0065;14'd5845:data <=32'h00A60036;14'd5846:data <=32'h00930011;
14'd5847:data <=32'h0077FFF7;14'd5848:data <=32'h005CFFEA;14'd5849:data <=32'h0043FFE7;
14'd5850:data <=32'h0030FFE8;14'd5851:data <=32'h0020FFED;14'd5852:data <=32'h0015FFF3;
14'd5853:data <=32'h000BFFF9;14'd5854:data <=32'h00010001;14'd5855:data <=32'hFFFA000B;
14'd5856:data <=32'hFFF40019;14'd5857:data <=32'hFFF3002A;14'd5858:data <=32'hFFF8003B;
14'd5859:data <=32'h0003004A;14'd5860:data <=32'h00110056;14'd5861:data <=32'h0024005D;
14'd5862:data <=32'h00380060;14'd5863:data <=32'h004C005F;14'd5864:data <=32'h005F005A;
14'd5865:data <=32'h00730052;14'd5866:data <=32'h00870047;14'd5867:data <=32'h009C0036;
14'd5868:data <=32'h00AE001F;14'd5869:data <=32'h00BD0001;14'd5870:data <=32'h00C4FFDD;
14'd5871:data <=32'h00C1FFB7;14'd5872:data <=32'h00B2FF90;14'd5873:data <=32'h0097FF70;
14'd5874:data <=32'h0074FF5A;14'd5875:data <=32'h004FFF4F;14'd5876:data <=32'h002AFF51;
14'd5877:data <=32'h000CFF5D;14'd5878:data <=32'hFFF7FF6F;14'd5879:data <=32'hFFECFF84;
14'd5880:data <=32'hFFE7FF94;14'd5881:data <=32'hFFEAFFA3;14'd5882:data <=32'hFFF1FFAC;
14'd5883:data <=32'hFFF9FFAF;14'd5884:data <=32'h0001FFAF;14'd5885:data <=32'h000AFFA7;
14'd5886:data <=32'h0011FF99;14'd5887:data <=32'h0013FF84;14'd5888:data <=32'hFFCAFF54;
14'd5889:data <=32'hFFB0FF47;14'd5890:data <=32'hFFA0FF52;14'd5891:data <=32'hFFDCFF7B;
14'd5892:data <=32'hFFB7FF2C;14'd5893:data <=32'hFF88FF2E;14'd5894:data <=32'hFF5BFF40;
14'd5895:data <=32'hFF32FF61;14'd5896:data <=32'hFF16FF88;14'd5897:data <=32'hFF06FFB6;
14'd5898:data <=32'hFF02FFE3;14'd5899:data <=32'hFF06000D;14'd5900:data <=32'hFF110032;
14'd5901:data <=32'hFF210055;14'd5902:data <=32'hFF360074;14'd5903:data <=32'hFF50008F;
14'd5904:data <=32'hFF6F00A3;14'd5905:data <=32'hFF9100AF;14'd5906:data <=32'hFFB400B3;
14'd5907:data <=32'hFFD500AE;14'd5908:data <=32'hFFF000A4;14'd5909:data <=32'h00030094;
14'd5910:data <=32'h00100087;14'd5911:data <=32'h0019007C;14'd5912:data <=32'h00210072;
14'd5913:data <=32'h002C006B;14'd5914:data <=32'h00360061;14'd5915:data <=32'h00410053;
14'd5916:data <=32'h004A0041;14'd5917:data <=32'h004D002B;14'd5918:data <=32'h00480014;
14'd5919:data <=32'h003AFFFF;14'd5920:data <=32'h0027FFF0;14'd5921:data <=32'h000EFFEB;
14'd5922:data <=32'hFFF5FFEF;14'd5923:data <=32'hFFE0FFFB;14'd5924:data <=32'hFFD0000F;
14'd5925:data <=32'hFFC60027;14'd5926:data <=32'hFFC40040;14'd5927:data <=32'hFFCA005B;
14'd5928:data <=32'hFFD50077;14'd5929:data <=32'hFFEB0090;14'd5930:data <=32'h000800A5;
14'd5931:data <=32'h002C00B1;14'd5932:data <=32'h005500B6;14'd5933:data <=32'h008400AC;
14'd5934:data <=32'h00AD0095;14'd5935:data <=32'h00D10071;14'd5936:data <=32'h00E70044;
14'd5937:data <=32'h00EF0014;14'd5938:data <=32'h00E9FFE6;14'd5939:data <=32'h00D7FFBD;
14'd5940:data <=32'h00BEFF9F;14'd5941:data <=32'h00A2FF8C;14'd5942:data <=32'h0087FF82;
14'd5943:data <=32'h0071FF7E;14'd5944:data <=32'h005FFF7D;14'd5945:data <=32'h0050FF7D;
14'd5946:data <=32'h0043FF7C;14'd5947:data <=32'h0038FF7D;14'd5948:data <=32'h0030FF7F;
14'd5949:data <=32'h002BFF7F;14'd5950:data <=32'h0027FF7D;14'd5951:data <=32'h0024FF78;
14'd5952:data <=32'h0044FFD2;14'd5953:data <=32'h005DFFB0;14'd5954:data <=32'h0054FF8B;
14'd5955:data <=32'hFFEDFF64;14'd5956:data <=32'hFFCFFF21;14'd5957:data <=32'hFFAAFF2C;
14'd5958:data <=32'hFF87FF42;14'd5959:data <=32'hFF6CFF5F;14'd5960:data <=32'hFF5CFF84;
14'd5961:data <=32'hFF58FFA8;14'd5962:data <=32'hFF5EFFC8;14'd5963:data <=32'hFF6BFFDF;
14'd5964:data <=32'hFF79FFEE;14'd5965:data <=32'hFF85FFF6;14'd5966:data <=32'hFF8EFFFA;
14'd5967:data <=32'hFF93FFFD;14'd5968:data <=32'hFF970000;14'd5969:data <=32'hFF9A0003;
14'd5970:data <=32'hFF990005;14'd5971:data <=32'hFF990008;14'd5972:data <=32'hFF95000B;
14'd5973:data <=32'hFF8E0011;14'd5974:data <=32'hFF87001C;14'd5975:data <=32'hFF81002F;
14'd5976:data <=32'hFF810046;14'd5977:data <=32'hFF8A0060;14'd5978:data <=32'hFF9D0077;
14'd5979:data <=32'hFFB90089;14'd5980:data <=32'hFFD9008F;14'd5981:data <=32'hFFFA008A;
14'd5982:data <=32'h0016007B;14'd5983:data <=32'h002B0063;14'd5984:data <=32'h00340047;
14'd5985:data <=32'h0033002D;14'd5986:data <=32'h002A0017;14'd5987:data <=32'h001B0007;
14'd5988:data <=32'h0008FFFD;14'd5989:data <=32'hFFF5FFFA;14'd5990:data <=32'hFFE1FFFE;
14'd5991:data <=32'hFFCE0007;14'd5992:data <=32'hFFBE0017;14'd5993:data <=32'hFFB2002C;
14'd5994:data <=32'hFFAC0047;14'd5995:data <=32'hFFAF0065;14'd5996:data <=32'hFFBC0081;
14'd5997:data <=32'hFFD4009C;14'd5998:data <=32'hFFF200AD;14'd5999:data <=32'h001400B6;
14'd6000:data <=32'h003600B4;14'd6001:data <=32'h005300AB;14'd6002:data <=32'h006C009D;
14'd6003:data <=32'h007F008D;14'd6004:data <=32'h0090007D;14'd6005:data <=32'h009E0071;
14'd6006:data <=32'h00AE0063;14'd6007:data <=32'h00C00053;14'd6008:data <=32'h00D4003F;
14'd6009:data <=32'h00E60023;14'd6010:data <=32'h00F30002;14'd6011:data <=32'h00F9FFDB;
14'd6012:data <=32'h00F7FFB3;14'd6013:data <=32'h00ECFF8B;14'd6014:data <=32'h00DAFF66;
14'd6015:data <=32'h00C3FF45;14'd6016:data <=32'h0023FFFC;14'd6017:data <=32'h004DFFFB;
14'd6018:data <=32'h0078FFD7;14'd6019:data <=32'h008CFF1A;14'd6020:data <=32'h0056FEC2;
14'd6021:data <=32'h0014FEC0;14'd6022:data <=32'hFFD3FED1;14'd6023:data <=32'hFF99FEF1;
14'd6024:data <=32'hFF70FF20;14'd6025:data <=32'hFF58FF55;14'd6026:data <=32'hFF52FF8A;
14'd6027:data <=32'hFF5CFFB6;14'd6028:data <=32'hFF6FFFD9;14'd6029:data <=32'hFF86FFEE;
14'd6030:data <=32'hFF9EFFFA;14'd6031:data <=32'hFFB4FFFD;14'd6032:data <=32'hFFC5FFFC;
14'd6033:data <=32'hFFD3FFF5;14'd6034:data <=32'hFFDDFFEB;14'd6035:data <=32'hFFE0FFDE;
14'd6036:data <=32'hFFDCFFCF;14'd6037:data <=32'hFFD2FFC2;14'd6038:data <=32'hFFC0FFB9;
14'd6039:data <=32'hFFAAFFBA;14'd6040:data <=32'hFF93FFC5;14'd6041:data <=32'hFF81FFD9;
14'd6042:data <=32'hFF78FFF3;14'd6043:data <=32'hFF78000E;14'd6044:data <=32'hFF820027;
14'd6045:data <=32'hFF92003A;14'd6046:data <=32'hFFA40044;14'd6047:data <=32'hFFB80048;
14'd6048:data <=32'hFFC60046;14'd6049:data <=32'hFFD00041;14'd6050:data <=32'hFFD8003C;
14'd6051:data <=32'hFFDD0039;14'd6052:data <=32'hFFE00035;14'd6053:data <=32'hFFE30032;
14'd6054:data <=32'hFFE6002F;14'd6055:data <=32'hFFE8002A;14'd6056:data <=32'hFFE70025;
14'd6057:data <=32'hFFE20021;14'd6058:data <=32'hFFDC0020;14'd6059:data <=32'hFFD50022;
14'd6060:data <=32'hFFCE0026;14'd6061:data <=32'hFFC9002F;14'd6062:data <=32'hFFC60037;
14'd6063:data <=32'hFFC40041;14'd6064:data <=32'hFFC4004A;14'd6065:data <=32'hFFC20054;
14'd6066:data <=32'hFFBE0061;14'd6067:data <=32'hFFBD0073;14'd6068:data <=32'hFFBD008B;
14'd6069:data <=32'hFFC600A9;14'd6070:data <=32'hFFDA00C9;14'd6071:data <=32'hFFFC00E8;
14'd6072:data <=32'h002900FF;14'd6073:data <=32'h00600108;14'd6074:data <=32'h009D0101;
14'd6075:data <=32'h00D800EA;14'd6076:data <=32'h010B00C4;14'd6077:data <=32'h01350092;
14'd6078:data <=32'h01520057;14'd6079:data <=32'h01630017;14'd6080:data <=32'h007C000C;
14'd6081:data <=32'h009B0009;14'd6082:data <=32'h00C90008;14'd6083:data <=32'h014CFFDA;
14'd6084:data <=32'h0137FF56;14'd6085:data <=32'h0105FF21;14'd6086:data <=32'h00CAFEFC;
14'd6087:data <=32'h008AFEEA;14'd6088:data <=32'h004CFEEC;14'd6089:data <=32'h0017FEFC;
14'd6090:data <=32'hFFEFFF18;14'd6091:data <=32'hFFD3FF35;14'd6092:data <=32'hFFC3FF51;
14'd6093:data <=32'hFFBAFF6A;14'd6094:data <=32'hFFB3FF7F;14'd6095:data <=32'hFFB0FF92;
14'd6096:data <=32'hFFAFFFA3;14'd6097:data <=32'hFFB0FFB3;14'd6098:data <=32'hFFB4FFC1;
14'd6099:data <=32'hFFBAFFCB;14'd6100:data <=32'hFFC2FFD2;14'd6101:data <=32'hFFC7FFD3;
14'd6102:data <=32'hFFCAFFD2;14'd6103:data <=32'hFFCAFFD2;14'd6104:data <=32'hFFC6FFD2;
14'd6105:data <=32'hFFC2FFD8;14'd6106:data <=32'hFFC0FFDF;14'd6107:data <=32'hFFC0FFE6;
14'd6108:data <=32'hFFC6FFED;14'd6109:data <=32'hFFCEFFEF;14'd6110:data <=32'hFFD4FFEB;
14'd6111:data <=32'hFFD6FFE3;14'd6112:data <=32'hFFD3FFDA;14'd6113:data <=32'hFFC9FFD2;
14'd6114:data <=32'hFFBAFFD1;14'd6115:data <=32'hFFABFFD6;14'd6116:data <=32'hFF9CFFE2;
14'd6117:data <=32'hFF94FFF3;14'd6118:data <=32'hFF910004;14'd6119:data <=32'hFF930016;
14'd6120:data <=32'hFF9A0025;14'd6121:data <=32'hFFA50030;14'd6122:data <=32'hFFB10038;
14'd6123:data <=32'hFFBC003B;14'd6124:data <=32'hFFC7003B;14'd6125:data <=32'hFFD0003A;
14'd6126:data <=32'hFFD90034;14'd6127:data <=32'hFFDD002B;14'd6128:data <=32'hFFDC0020;
14'd6129:data <=32'hFFD40016;14'd6130:data <=32'hFFC6000D;14'd6131:data <=32'hFFB0000D;
14'd6132:data <=32'hFF950017;14'd6133:data <=32'hFF7D0030;14'd6134:data <=32'hFF6C0054;
14'd6135:data <=32'hFF690081;14'd6136:data <=32'hFF7500B1;14'd6137:data <=32'hFF9100DF;
14'd6138:data <=32'hFFBC0104;14'd6139:data <=32'hFFF0011B;14'd6140:data <=32'h00290126;
14'd6141:data <=32'h00630121;14'd6142:data <=32'h009A0112;14'd6143:data <=32'h00CD00F5;
14'd6144:data <=32'h008100D5;14'd6145:data <=32'h00BC00D7;14'd6146:data <=32'h00E500D1;
14'd6147:data <=32'h00D400CE;14'd6148:data <=32'h00F40061;14'd6149:data <=32'h00F90037;
14'd6150:data <=32'h00F5000F;14'd6151:data <=32'h00E8FFED;14'd6152:data <=32'h00D7FFD3;
14'd6153:data <=32'h00C8FFC0;14'd6154:data <=32'h00BCFFB1;14'd6155:data <=32'h00B2FFA3;
14'd6156:data <=32'h00A9FF91;14'd6157:data <=32'h009FFF7D;14'd6158:data <=32'h008FFF65;
14'd6159:data <=32'h0077FF50;14'd6160:data <=32'h0058FF3E;14'd6161:data <=32'h0035FF36;
14'd6162:data <=32'h0012FF36;14'd6163:data <=32'hFFF0FF40;14'd6164:data <=32'hFFD3FF4E;
14'd6165:data <=32'hFFBAFF62;14'd6166:data <=32'hFFA9FF79;14'd6167:data <=32'hFF9AFF93;
14'd6168:data <=32'hFF91FFAE;14'd6169:data <=32'hFF91FFCC;14'd6170:data <=32'hFF97FFE8;
14'd6171:data <=32'hFFA70002;14'd6172:data <=32'hFFBE0016;14'd6173:data <=32'hFFDC0020;
14'd6174:data <=32'hFFFA001C;14'd6175:data <=32'h0014000D;14'd6176:data <=32'h0025FFF5;
14'd6177:data <=32'h002BFFD8;14'd6178:data <=32'h0024FFBC;14'd6179:data <=32'h0014FFA4;
14'd6180:data <=32'hFFFDFF95;14'd6181:data <=32'hFFE4FF91;14'd6182:data <=32'hFFCBFF92;
14'd6183:data <=32'hFFB6FF9B;14'd6184:data <=32'hFFA5FFA6;14'd6185:data <=32'hFF96FFB4;
14'd6186:data <=32'hFF8DFFC4;14'd6187:data <=32'hFF86FFD4;14'd6188:data <=32'hFF83FFE4;
14'd6189:data <=32'hFF82FFF5;14'd6190:data <=32'hFF860003;14'd6191:data <=32'hFF8C000E;
14'd6192:data <=32'hFF940015;14'd6193:data <=32'hFF990018;14'd6194:data <=32'hFF9A0018;
14'd6195:data <=32'hFF950017;14'd6196:data <=32'hFF8B0019;14'd6197:data <=32'hFF7E0024;
14'd6198:data <=32'hFF720036;14'd6199:data <=32'hFF6C0051;14'd6200:data <=32'hFF6D006F;
14'd6201:data <=32'hFF79008F;14'd6202:data <=32'hFF8F00AB;14'd6203:data <=32'hFFAB00BE;
14'd6204:data <=32'hFFCB00CB;14'd6205:data <=32'hFFEA00D0;14'd6206:data <=32'h000600CF;
14'd6207:data <=32'h002100CA;14'd6208:data <=32'hFF930119;14'd6209:data <=32'hFFCE0150;
14'd6210:data <=32'h0011015A;14'd6211:data <=32'h002600BF;14'd6212:data <=32'h003D0075;
14'd6213:data <=32'h003E006F;14'd6214:data <=32'h003F006E;14'd6215:data <=32'h00410070;
14'd6216:data <=32'h00470077;14'd6217:data <=32'h00530081;14'd6218:data <=32'h0068008A;
14'd6219:data <=32'h0087008B;14'd6220:data <=32'h00AC0081;14'd6221:data <=32'h00D00069;
14'd6222:data <=32'h00EE0044;14'd6223:data <=32'h01000015;14'd6224:data <=32'h0104FFE0;
14'd6225:data <=32'h00F8FFAD;14'd6226:data <=32'h00DFFF7F;14'd6227:data <=32'h00BDFF5A;
14'd6228:data <=32'h0095FF41;14'd6229:data <=32'h006AFF30;14'd6230:data <=32'h003DFF2A;
14'd6231:data <=32'h0012FF2E;14'd6232:data <=32'hFFE8FF3C;14'd6233:data <=32'hFFC2FF54;
14'd6234:data <=32'hFFA6FF77;14'd6235:data <=32'hFF97FF9E;14'd6236:data <=32'hFF95FFC8;
14'd6237:data <=32'hFFA0FFED;14'd6238:data <=32'hFFB7000A;14'd6239:data <=32'hFFD4001B;
14'd6240:data <=32'hFFF30021;14'd6241:data <=32'h000F001B;14'd6242:data <=32'h0023000C;
14'd6243:data <=32'h0032FFFB;14'd6244:data <=32'h0037FFE7;14'd6245:data <=32'h003AFFD5;
14'd6246:data <=32'h0039FFC6;14'd6247:data <=32'h0036FFB5;14'd6248:data <=32'h0031FFA6;
14'd6249:data <=32'h0029FF95;14'd6250:data <=32'h001DFF84;14'd6251:data <=32'h000CFF74;
14'd6252:data <=32'hFFF5FF67;14'd6253:data <=32'hFFDAFF5F;14'd6254:data <=32'hFFBEFF5E;
14'd6255:data <=32'hFFA2FF62;14'd6256:data <=32'hFF87FF6A;14'd6257:data <=32'hFF6DFF78;
14'd6258:data <=32'hFF54FF89;14'd6259:data <=32'hFF3CFF9F;14'd6260:data <=32'hFF26FFBA;
14'd6261:data <=32'hFF12FFDB;14'd6262:data <=32'hFF060004;14'd6263:data <=32'hFF030032;
14'd6264:data <=32'hFF0D0063;14'd6265:data <=32'hFF240090;14'd6266:data <=32'hFF4800B5;
14'd6267:data <=32'hFF7400CE;14'd6268:data <=32'hFFA300D7;14'd6269:data <=32'hFFCE00D4;
14'd6270:data <=32'hFFF200C5;14'd6271:data <=32'h000C00B1;14'd6272:data <=32'hFF29006B;
14'd6273:data <=32'hFF2B00AD;14'd6274:data <=32'hFF5A00E9;14'd6275:data <=32'h000900B3;
14'd6276:data <=32'h001E005E;14'd6277:data <=32'h00140050;14'd6278:data <=32'h00070048;
14'd6279:data <=32'hFFFA004A;14'd6280:data <=32'hFFEC0054;14'd6281:data <=32'hFFE40068;
14'd6282:data <=32'hFFE80082;14'd6283:data <=32'hFFF9009C;14'd6284:data <=32'h001600B2;
14'd6285:data <=32'h003D00BC;14'd6286:data <=32'h006700B7;14'd6287:data <=32'h008E00A6;
14'd6288:data <=32'h00AF0089;14'd6289:data <=32'h00C50064;14'd6290:data <=32'h00D0003E;
14'd6291:data <=32'h00D30019;14'd6292:data <=32'h00CEFFF5;14'd6293:data <=32'h00C3FFD4;
14'd6294:data <=32'h00B2FFB7;14'd6295:data <=32'h009DFF9F;14'd6296:data <=32'h0082FF8B;
14'd6297:data <=32'h0064FF7E;14'd6298:data <=32'h0044FF7A;14'd6299:data <=32'h0025FF7F;
14'd6300:data <=32'h000CFF8C;14'd6301:data <=32'hFFF9FF9E;14'd6302:data <=32'hFFF0FFB2;
14'd6303:data <=32'hFFEDFFC4;14'd6304:data <=32'hFFEDFFD3;14'd6305:data <=32'hFFF1FFDE;
14'd6306:data <=32'hFFF5FFE5;14'd6307:data <=32'hFFF7FFEE;14'd6308:data <=32'hFFFCFFF8;
14'd6309:data <=32'h00030002;14'd6310:data <=32'h000E000C;14'd6311:data <=32'h00200013;
14'd6312:data <=32'h00360014;14'd6313:data <=32'h0050000C;14'd6314:data <=32'h0069FFFC;
14'd6315:data <=32'h007CFFE0;14'd6316:data <=32'h0088FFBE;14'd6317:data <=32'h0088FF97;
14'd6318:data <=32'h007FFF6F;14'd6319:data <=32'h0069FF49;14'd6320:data <=32'h004BFF28;
14'd6321:data <=32'h0025FF0D;14'd6322:data <=32'hFFF7FEF9;14'd6323:data <=32'hFFC3FEF1;
14'd6324:data <=32'hFF8AFEF4;14'd6325:data <=32'hFF50FF04;14'd6326:data <=32'hFF19FF25;
14'd6327:data <=32'hFEEBFF55;14'd6328:data <=32'hFECBFF92;14'd6329:data <=32'hFEBEFFD5;
14'd6330:data <=32'hFEC30018;14'd6331:data <=32'hFEDB0054;14'd6332:data <=32'hFF000083;
14'd6333:data <=32'hFF2C00A4;14'd6334:data <=32'hFF5A00B5;14'd6335:data <=32'hFF8300BA;
14'd6336:data <=32'hFF64002E;14'd6337:data <=32'hFF560049;14'd6338:data <=32'hFF4F007B;
14'd6339:data <=32'hFF7300CF;14'd6340:data <=32'hFFA00090;14'd6341:data <=32'hFFB10090;
14'd6342:data <=32'hFFBE008D;14'd6343:data <=32'hFFCA008C;14'd6344:data <=32'hFFD1008B;
14'd6345:data <=32'hFFD70090;14'd6346:data <=32'hFFE00098;14'd6347:data <=32'hFFEE00A2;
14'd6348:data <=32'h000300AB;14'd6349:data <=32'h001D00AD;14'd6350:data <=32'h003A00A6;
14'd6351:data <=32'h00540098;14'd6352:data <=32'h00670081;14'd6353:data <=32'h00710067;
14'd6354:data <=32'h0073004F;14'd6355:data <=32'h006F003A;14'd6356:data <=32'h0068002C;
14'd6357:data <=32'h00610024;14'd6358:data <=32'h005D001D;14'd6359:data <=32'h005A0018;
14'd6360:data <=32'h00590014;14'd6361:data <=32'h0057000E;14'd6362:data <=32'h00550009;
14'd6363:data <=32'h00530004;14'd6364:data <=32'h00500000;14'd6365:data <=32'h0050FFFD;
14'd6366:data <=32'h0053FFFA;14'd6367:data <=32'h0054FFF3;14'd6368:data <=32'h0055FFE8;
14'd6369:data <=32'h0050FFDC;14'd6370:data <=32'h0047FFCF;14'd6371:data <=32'h0038FFC7;
14'd6372:data <=32'h0025FFC5;14'd6373:data <=32'h0012FFCB;14'd6374:data <=32'h0003FFDA;
14'd6375:data <=32'hFFFDFFF0;14'd6376:data <=32'h00000008;14'd6377:data <=32'h000F001B;
14'd6378:data <=32'h00270029;14'd6379:data <=32'h0044002D;14'd6380:data <=32'h00620026;
14'd6381:data <=32'h007D0015;14'd6382:data <=32'h0094FFFB;14'd6383:data <=32'h00A3FFDB;
14'd6384:data <=32'h00AAFFB7;14'd6385:data <=32'h00A9FF8E;14'd6386:data <=32'h009EFF66;
14'd6387:data <=32'h0089FF3E;14'd6388:data <=32'h0069FF1B;14'd6389:data <=32'h003FFEFD;
14'd6390:data <=32'h000CFEEC;14'd6391:data <=32'hFFD4FEE8;14'd6392:data <=32'hFF9EFEF4;
14'd6393:data <=32'hFF6FFF0D;14'd6394:data <=32'hFF49FF30;14'd6395:data <=32'hFF31FF58;
14'd6396:data <=32'hFF23FF7F;14'd6397:data <=32'hFF1EFFA1;14'd6398:data <=32'hFF1EFFBF;
14'd6399:data <=32'hFF1EFFD8;14'd6400:data <=32'hFF290010;14'd6401:data <=32'hFF27002B;
14'd6402:data <=32'hFF200038;14'd6403:data <=32'hFEE8FFF3;14'd6404:data <=32'hFEF4FFDA;
14'd6405:data <=32'hFEED0005;14'd6406:data <=32'hFEEF0030;14'd6407:data <=32'hFEF9005D;
14'd6408:data <=32'hFF0B0086;14'd6409:data <=32'hFF2300AD;14'd6410:data <=32'hFF4300D0;
14'd6411:data <=32'hFF6B00ED;14'd6412:data <=32'hFF9C0102;14'd6413:data <=32'hFFD3010A;
14'd6414:data <=32'h000B0102;14'd6415:data <=32'h003D00EB;14'd6416:data <=32'h006600C7;
14'd6417:data <=32'h007F009A;14'd6418:data <=32'h0088006C;14'd6419:data <=32'h00810042;
14'd6420:data <=32'h00710021;14'd6421:data <=32'h005A000C;14'd6422:data <=32'h00420000;
14'd6423:data <=32'h002DFFFD;14'd6424:data <=32'h001A0001;14'd6425:data <=32'h000C0009;
14'd6426:data <=32'h00020013;14'd6427:data <=32'hFFFB0021;14'd6428:data <=32'hFFFB0031;
14'd6429:data <=32'h00010040;14'd6430:data <=32'h000D004E;14'd6431:data <=32'h001F0055;
14'd6432:data <=32'h00330055;14'd6433:data <=32'h0047004D;14'd6434:data <=32'h0055003F;
14'd6435:data <=32'h005C002D;14'd6436:data <=32'h005C001C;14'd6437:data <=32'h0055000D;
14'd6438:data <=32'h004B0006;14'd6439:data <=32'h00420005;14'd6440:data <=32'h003C000A;
14'd6441:data <=32'h003B0011;14'd6442:data <=32'h00420016;14'd6443:data <=32'h004B0019;
14'd6444:data <=32'h00580017;14'd6445:data <=32'h00630010;14'd6446:data <=32'h006B0006;
14'd6447:data <=32'h0074FFF9;14'd6448:data <=32'h0078FFED;14'd6449:data <=32'h007CFFDF;
14'd6450:data <=32'h007EFFD0;14'd6451:data <=32'h007FFFBF;14'd6452:data <=32'h007DFFAD;
14'd6453:data <=32'h0077FF9A;14'd6454:data <=32'h006CFF87;14'd6455:data <=32'h005DFF77;
14'd6456:data <=32'h004DFF6C;14'd6457:data <=32'h003CFF65;14'd6458:data <=32'h002EFF60;
14'd6459:data <=32'h0024FF5C;14'd6460:data <=32'h001BFF54;14'd6461:data <=32'h0012FF49;
14'd6462:data <=32'h0002FF37;14'd6463:data <=32'hFFEAFF25;14'd6464:data <=32'hFF4EFF55;
14'd6465:data <=32'hFF33FF69;14'd6466:data <=32'hFF33FF7B;14'd6467:data <=32'hFF97FF1A;
14'd6468:data <=32'hFF79FEE3;14'd6469:data <=32'hFF3FFEF9;14'd6470:data <=32'hFF0BFF1D;
14'd6471:data <=32'hFEDFFF4D;14'd6472:data <=32'hFEC0FF85;14'd6473:data <=32'hFEADFFC3;
14'd6474:data <=32'hFEA70006;14'd6475:data <=32'hFEB1004A;14'd6476:data <=32'hFECE008C;
14'd6477:data <=32'hFEF900C3;14'd6478:data <=32'hFF3400EC;14'd6479:data <=32'hFF750103;
14'd6480:data <=32'hFFB60103;14'd6481:data <=32'hFFEF00F2;14'd6482:data <=32'h001D00D5;
14'd6483:data <=32'h003B00B1;14'd6484:data <=32'h004D008B;14'd6485:data <=32'h00530069;
14'd6486:data <=32'h0050004B;14'd6487:data <=32'h00490033;14'd6488:data <=32'h0040001F;
14'd6489:data <=32'h00330010;14'd6490:data <=32'h00230005;14'd6491:data <=32'h0011FFFE;
14'd6492:data <=32'hFFFFFFFF;14'd6493:data <=32'hFFEF0005;14'd6494:data <=32'hFFE30011;
14'd6495:data <=32'hFFDB0020;14'd6496:data <=32'hFFDB0030;14'd6497:data <=32'hFFDF003E;
14'd6498:data <=32'hFFE60048;14'd6499:data <=32'hFFEE0050;14'd6500:data <=32'hFFF40056;
14'd6501:data <=32'hFFFB005D;14'd6502:data <=32'h00020065;14'd6503:data <=32'h000C006E;
14'd6504:data <=32'h001C007A;14'd6505:data <=32'h00300081;14'd6506:data <=32'h004A0084;
14'd6507:data <=32'h0066007D;14'd6508:data <=32'h0082006E;14'd6509:data <=32'h00970056;
14'd6510:data <=32'h00A60039;14'd6511:data <=32'h00AB001B;14'd6512:data <=32'h00A8FFFD;
14'd6513:data <=32'h009EFFE4;14'd6514:data <=32'h008FFFD1;14'd6515:data <=32'h0080FFC4;
14'd6516:data <=32'h006FFFBA;14'd6517:data <=32'h0060FFB6;14'd6518:data <=32'h0051FFB6;
14'd6519:data <=32'h0045FFBA;14'd6520:data <=32'h003CFFC2;14'd6521:data <=32'h003AFFCD;
14'd6522:data <=32'h003FFFD7;14'd6523:data <=32'h004EFFDF;14'd6524:data <=32'h0063FFDE;
14'd6525:data <=32'h007CFFCF;14'd6526:data <=32'h0091FFB3;14'd6527:data <=32'h009CFF8B;
14'd6528:data <=32'h0045FF46;14'd6529:data <=32'h0032FF27;14'd6530:data <=32'h001DFF28;
14'd6531:data <=32'h0053FF5C;14'd6532:data <=32'h004AFF01;14'd6533:data <=32'h001BFEF1;
14'd6534:data <=32'hFFEAFEE9;14'd6535:data <=32'hFFB8FEEF;14'd6536:data <=32'hFF89FEFD;
14'd6537:data <=32'hFF5CFF14;14'd6538:data <=32'hFF35FF36;14'd6539:data <=32'hFF14FF60;
14'd6540:data <=32'hFEFFFF91;14'd6541:data <=32'hFEF9FFC6;14'd6542:data <=32'hFF00FFF9;
14'd6543:data <=32'hFF130024;14'd6544:data <=32'hFF2E0046;14'd6545:data <=32'hFF4D005C;
14'd6546:data <=32'hFF6A0068;14'd6547:data <=32'hFF82006D;14'd6548:data <=32'hFF960070;
14'd6549:data <=32'hFFA80073;14'd6550:data <=32'hFFB80076;14'd6551:data <=32'hFFCC0078;
14'd6552:data <=32'hFFDF0078;14'd6553:data <=32'hFFF40072;14'd6554:data <=32'h00070066;
14'd6555:data <=32'h00150056;14'd6556:data <=32'h001E0043;14'd6557:data <=32'h00200030;
14'd6558:data <=32'h001D001E;14'd6559:data <=32'h0014000F;14'd6560:data <=32'h000A0003;
14'd6561:data <=32'hFFFCFFFB;14'd6562:data <=32'hFFEDFFF5;14'd6563:data <=32'hFFDBFFF4;
14'd6564:data <=32'hFFC6FFF9;14'd6565:data <=32'hFFB10005;14'd6566:data <=32'hFF9E0019;
14'd6567:data <=32'hFF910036;14'd6568:data <=32'hFF8E005A;14'd6569:data <=32'hFF970081;
14'd6570:data <=32'hFFAE00A5;14'd6571:data <=32'hFFD000C1;14'd6572:data <=32'hFFFB00D0;
14'd6573:data <=32'h002800D4;14'd6574:data <=32'h005300C8;14'd6575:data <=32'h007800B3;
14'd6576:data <=32'h00930097;14'd6577:data <=32'h00A50078;14'd6578:data <=32'h00AF0058;
14'd6579:data <=32'h00B2003A;14'd6580:data <=32'h00AF001F;14'd6581:data <=32'h00A80006;
14'd6582:data <=32'h009CFFF2;14'd6583:data <=32'h008DFFE3;14'd6584:data <=32'h007DFFDA;
14'd6585:data <=32'h006EFFD9;14'd6586:data <=32'h0064FFDF;14'd6587:data <=32'h0064FFE6;
14'd6588:data <=32'h006AFFED;14'd6589:data <=32'h0079FFED;14'd6590:data <=32'h008BFFE4;
14'd6591:data <=32'h009CFFD1;14'd6592:data <=32'h008A0013;14'd6593:data <=32'h00B1FFF4;
14'd6594:data <=32'h00B7FFCB;14'd6595:data <=32'h0064FF8F;14'd6596:data <=32'h0068FF41;
14'd6597:data <=32'h0046FF38;14'd6598:data <=32'h0026FF39;14'd6599:data <=32'h000BFF40;
14'd6600:data <=32'hFFF3FF48;14'd6601:data <=32'hFFE0FF53;14'd6602:data <=32'hFFCEFF5E;
14'd6603:data <=32'hFFBEFF6B;14'd6604:data <=32'hFFB3FF7B;14'd6605:data <=32'hFFABFF8B;
14'd6606:data <=32'hFFA6FF9B;14'd6607:data <=32'hFFA8FFA7;14'd6608:data <=32'hFFAAFFAE;
14'd6609:data <=32'hFFABFFAF;14'd6610:data <=32'hFFA7FFAD;14'd6611:data <=32'hFF9CFFAC;
14'd6612:data <=32'hFF8BFFAE;14'd6613:data <=32'hFF78FFBA;14'd6614:data <=32'hFF65FFCF;
14'd6615:data <=32'hFF5AFFEB;14'd6616:data <=32'hFF59000C;14'd6617:data <=32'hFF61002C;
14'd6618:data <=32'hFF730046;14'd6619:data <=32'hFF8D005A;14'd6620:data <=32'hFFA90065;
14'd6621:data <=32'hFFC40068;14'd6622:data <=32'hFFDE0063;14'd6623:data <=32'hFFF4005A;
14'd6624:data <=32'h0006004A;14'd6625:data <=32'h00140036;14'd6626:data <=32'h0019001F;
14'd6627:data <=32'h00180006;14'd6628:data <=32'h000CFFEE;14'd6629:data <=32'hFFF7FFDB;
14'd6630:data <=32'hFFDCFFD1;14'd6631:data <=32'hFFBCFFD1;14'd6632:data <=32'hFF9CFFDE;
14'd6633:data <=32'hFF83FFF6;14'd6634:data <=32'hFF730015;14'd6635:data <=32'hFF6F003B;
14'd6636:data <=32'hFF76005D;14'd6637:data <=32'hFF86007C;14'd6638:data <=32'hFF9B0092;
14'd6639:data <=32'hFFB300A3;14'd6640:data <=32'hFFC900AD;14'd6641:data <=32'hFFE100B6;
14'd6642:data <=32'hFFF700BC;14'd6643:data <=32'h000E00C0;14'd6644:data <=32'h002800C1;
14'd6645:data <=32'h004300BF;14'd6646:data <=32'h005D00B9;14'd6647:data <=32'h007700AF;
14'd6648:data <=32'h008E009E;14'd6649:data <=32'h00A3008D;14'd6650:data <=32'h00B5007A;
14'd6651:data <=32'h00C50067;14'd6652:data <=32'h00D70051;14'd6653:data <=32'h00E80037;
14'd6654:data <=32'h00F60016;14'd6655:data <=32'h0100FFED;14'd6656:data <=32'h002A0050;
14'd6657:data <=32'h005C005E;14'd6658:data <=32'h00940048;14'd6659:data <=32'h00DEFF97;
14'd6660:data <=32'h00D4FF37;14'd6661:data <=32'h009EFF20;14'd6662:data <=32'h0068FF1B;
14'd6663:data <=32'h0036FF24;14'd6664:data <=32'h000FFF36;14'd6665:data <=32'hFFF3FF4C;
14'd6666:data <=32'hFFDEFF67;14'd6667:data <=32'hFFD1FF81;14'd6668:data <=32'hFFCDFF9C;
14'd6669:data <=32'hFFD1FFB4;14'd6670:data <=32'hFFDAFFC7;14'd6671:data <=32'hFFEBFFD3;
14'd6672:data <=32'hFFFFFFD5;14'd6673:data <=32'h0011FFCC;14'd6674:data <=32'h001CFFBB;
14'd6675:data <=32'h001CFFA3;14'd6676:data <=32'h0011FF8B;14'd6677:data <=32'hFFFAFF7A;
14'd6678:data <=32'hFFDDFF71;14'd6679:data <=32'hFFBDFF75;14'd6680:data <=32'hFFA1FF83;
14'd6681:data <=32'hFF8CFF99;14'd6682:data <=32'hFF81FFB3;14'd6683:data <=32'hFF7BFFCC;
14'd6684:data <=32'hFF7DFFE4;14'd6685:data <=32'hFF83FFF9;14'd6686:data <=32'hFF8C000B;
14'd6687:data <=32'hFF980019;14'd6688:data <=32'hFFA60024;14'd6689:data <=32'hFFB6002B;
14'd6690:data <=32'hFFC7002D;14'd6691:data <=32'hFFD80029;14'd6692:data <=32'hFFE60020;
14'd6693:data <=32'hFFEE0012;14'd6694:data <=32'hFFEE0002;14'd6695:data <=32'hFFE9FFF6;
14'd6696:data <=32'hFFDEFFEC;14'd6697:data <=32'hFFD1FFE8;14'd6698:data <=32'hFFC5FFE9;
14'd6699:data <=32'hFFBAFFEE;14'd6700:data <=32'hFFB2FFF3;14'd6701:data <=32'hFFACFFF8;
14'd6702:data <=32'hFFA4FFFB;14'd6703:data <=32'hFF9BFFFE;14'd6704:data <=32'hFF8C0004;
14'd6705:data <=32'hFF7B000F;14'd6706:data <=32'hFF690024;14'd6707:data <=32'hFF590041;
14'd6708:data <=32'hFF520065;14'd6709:data <=32'hFF55008E;14'd6710:data <=32'hFF6400B9;
14'd6711:data <=32'hFF7E00E2;14'd6712:data <=32'hFFA10103;14'd6713:data <=32'hFFCD011E;
14'd6714:data <=32'hFFFF0131;14'd6715:data <=32'h0037013A;14'd6716:data <=32'h00730138;
14'd6717:data <=32'h00B10128;14'd6718:data <=32'h00EE0108;14'd6719:data <=32'h012400D8;
14'd6720:data <=32'h00440064;14'd6721:data <=32'h00630076;14'd6722:data <=32'h00940088;
14'd6723:data <=32'h012E0082;14'd6724:data <=32'h014E0003;14'd6725:data <=32'h0133FFC7;
14'd6726:data <=32'h010EFF98;14'd6727:data <=32'h00E3FF77;14'd6728:data <=32'h00B9FF64;
14'd6729:data <=32'h0091FF5B;14'd6730:data <=32'h006CFF59;14'd6731:data <=32'h004BFF5D;
14'd6732:data <=32'h0030FF68;14'd6733:data <=32'h0019FF76;14'd6734:data <=32'h0009FF8A;
14'd6735:data <=32'h0001FF9E;14'd6736:data <=32'h0004FFAD;14'd6737:data <=32'h0009FFB9;
14'd6738:data <=32'h0011FFBC;14'd6739:data <=32'h0018FFB7;14'd6740:data <=32'h0019FFAE;
14'd6741:data <=32'h0013FFA5;14'd6742:data <=32'h0008FF9E;14'd6743:data <=32'hFFF9FF9E;
14'd6744:data <=32'hFFEDFFA4;14'd6745:data <=32'hFFE5FFAB;14'd6746:data <=32'hFFE1FFB4;
14'd6747:data <=32'hFFE1FFBB;14'd6748:data <=32'hFFE3FFBF;14'd6749:data <=32'hFFE5FFBF;
14'd6750:data <=32'hFFE3FFBD;14'd6751:data <=32'hFFDEFFBA;14'd6752:data <=32'hFFD7FFBA;
14'd6753:data <=32'hFFCFFFBB;14'd6754:data <=32'hFFC8FFC0;14'd6755:data <=32'hFFC2FFC6;
14'd6756:data <=32'hFFBDFFCB;14'd6757:data <=32'hFFBAFFD1;14'd6758:data <=32'hFFB6FFD8;
14'd6759:data <=32'hFFB3FFDF;14'd6760:data <=32'hFFB0FFE7;14'd6761:data <=32'hFFB0FFF1;
14'd6762:data <=32'hFFB4FFFC;14'd6763:data <=32'hFFBD0005;14'd6764:data <=32'hFFC90008;
14'd6765:data <=32'hFFD60005;14'd6766:data <=32'hFFE1FFFA;14'd6767:data <=32'hFFE5FFE7;
14'd6768:data <=32'hFFDFFFD2;14'd6769:data <=32'hFFCEFFBD;14'd6770:data <=32'hFFB0FFB0;
14'd6771:data <=32'hFF8CFFAE;14'd6772:data <=32'hFF66FFBA;14'd6773:data <=32'hFF41FFD2;
14'd6774:data <=32'hFF25FFF8;14'd6775:data <=32'hFF130026;14'd6776:data <=32'hFF0C0057;
14'd6777:data <=32'hFF12008B;14'd6778:data <=32'hFF2300C0;14'd6779:data <=32'hFF4000F2;
14'd6780:data <=32'hFF6A011F;14'd6781:data <=32'hFFA00143;14'd6782:data <=32'hFFE10159;
14'd6783:data <=32'h0028015E;14'd6784:data <=32'hFFFA00FC;14'd6785:data <=32'h002E0117;
14'd6786:data <=32'h00520126;14'd6787:data <=32'h004F012F;14'd6788:data <=32'h009800D8;
14'd6789:data <=32'h00AB00B8;14'd6790:data <=32'h00B80099;14'd6791:data <=32'h00BF007E;
14'd6792:data <=32'h00C50067;14'd6793:data <=32'h00CD004F;14'd6794:data <=32'h00D30035;
14'd6795:data <=32'h00D60019;14'd6796:data <=32'h00D5FFFC;14'd6797:data <=32'h00CCFFDF;
14'd6798:data <=32'h00C1FFC5;14'd6799:data <=32'h00B1FFAF;14'd6800:data <=32'h00A1FF9C;
14'd6801:data <=32'h008EFF8C;14'd6802:data <=32'h007AFF7E;14'd6803:data <=32'h0065FF70;
14'd6804:data <=32'h0049FF67;14'd6805:data <=32'h002BFF62;14'd6806:data <=32'h000AFF67;
14'd6807:data <=32'hFFECFF75;14'd6808:data <=32'hFFD4FF8E;14'd6809:data <=32'hFFC6FFAB;
14'd6810:data <=32'hFFC4FFCB;14'd6811:data <=32'hFFCEFFE6;14'd6812:data <=32'hFFE1FFF9;
14'd6813:data <=32'hFFF90004;14'd6814:data <=32'h00100002;14'd6815:data <=32'h0022FFF9;
14'd6816:data <=32'h002FFFEA;14'd6817:data <=32'h0036FFD9;14'd6818:data <=32'h0037FFC6;
14'd6819:data <=32'h0032FFB6;14'd6820:data <=32'h002AFFA4;14'd6821:data <=32'h001DFF97;
14'd6822:data <=32'h000CFF8C;14'd6823:data <=32'hFFF8FF87;14'd6824:data <=32'hFFE2FF86;
14'd6825:data <=32'hFFCDFF8D;14'd6826:data <=32'hFFBDFF9A;14'd6827:data <=32'hFFB2FFAA;
14'd6828:data <=32'hFFAFFFBC;14'd6829:data <=32'hFFB3FFCB;14'd6830:data <=32'hFFBCFFD3;
14'd6831:data <=32'hFFC5FFD3;14'd6832:data <=32'hFFCBFFCC;14'd6833:data <=32'hFFCAFFC0;
14'd6834:data <=32'hFFC0FFB3;14'd6835:data <=32'hFFADFFAB;14'd6836:data <=32'hFF95FFA9;
14'd6837:data <=32'hFF7CFFB0;14'd6838:data <=32'hFF65FFC0;14'd6839:data <=32'hFF51FFD5;
14'd6840:data <=32'hFF43FFEF;14'd6841:data <=32'hFF39000C;14'd6842:data <=32'hFF350029;
14'd6843:data <=32'hFF35004A;14'd6844:data <=32'hFF3C006A;14'd6845:data <=32'hFF48008B;
14'd6846:data <=32'hFF5E00AB;14'd6847:data <=32'hFF7B00C6;14'd6848:data <=32'hFF0700D2;
14'd6849:data <=32'hFF29011C;14'd6850:data <=32'hFF5C013B;14'd6851:data <=32'hFF9700B9;
14'd6852:data <=32'hFFC70083;14'd6853:data <=32'hFFC70087;14'd6854:data <=32'hFFC70093;
14'd6855:data <=32'hFFCB00A4;14'd6856:data <=32'hFFD700BC;14'd6857:data <=32'hFFEF00D2;
14'd6858:data <=32'h001300E4;14'd6859:data <=32'h003D00EA;14'd6860:data <=32'h006900E5;
14'd6861:data <=32'h009500D4;14'd6862:data <=32'h00B900B9;14'd6863:data <=32'h00D90097;
14'd6864:data <=32'h00F0006E;14'd6865:data <=32'h01000040;14'd6866:data <=32'h01050011;
14'd6867:data <=32'h00FFFFDC;14'd6868:data <=32'h00EDFFAC;14'd6869:data <=32'h00CDFF80;
14'd6870:data <=32'h00A1FF60;14'd6871:data <=32'h006EFF4E;14'd6872:data <=32'h003BFF4D;
14'd6873:data <=32'h000DFF5C;14'd6874:data <=32'hFFE8FF78;14'd6875:data <=32'hFFD1FF9B;
14'd6876:data <=32'hFFC9FFBD;14'd6877:data <=32'hFFCCFFDF;14'd6878:data <=32'hFFD8FFF8;
14'd6879:data <=32'hFFE9000B;14'd6880:data <=32'hFFFC0016;14'd6881:data <=32'h0010001C;
14'd6882:data <=32'h0024001B;14'd6883:data <=32'h00360017;14'd6884:data <=32'h0048000E;
14'd6885:data <=32'h00580000;14'd6886:data <=32'h0063FFED;14'd6887:data <=32'h0069FFD7;
14'd6888:data <=32'h0068FFBE;14'd6889:data <=32'h0062FFA9;14'd6890:data <=32'h0056FF96;
14'd6891:data <=32'h0049FF86;14'd6892:data <=32'h003AFF7B;14'd6893:data <=32'h002BFF72;
14'd6894:data <=32'h001CFF67;14'd6895:data <=32'h000EFF5D;14'd6896:data <=32'hFFFCFF52;
14'd6897:data <=32'hFFE4FF48;14'd6898:data <=32'hFFC4FF41;14'd6899:data <=32'hFFA2FF42;
14'd6900:data <=32'hFF7DFF4E;14'd6901:data <=32'hFF5BFF65;14'd6902:data <=32'hFF3FFF85;
14'd6903:data <=32'hFF2CFFA9;14'd6904:data <=32'hFF27FFD1;14'd6905:data <=32'hFF29FFF7;
14'd6906:data <=32'hFF340016;14'd6907:data <=32'hFF430031;14'd6908:data <=32'hFF550046;
14'd6909:data <=32'hFF690057;14'd6910:data <=32'hFF7E0062;14'd6911:data <=32'hFF930068;
14'd6912:data <=32'hFEEBFFE8;14'd6913:data <=32'hFED20028;14'd6914:data <=32'hFEE7006D;
14'd6915:data <=32'hFF9E006A;14'd6916:data <=32'hFFC80024;14'd6917:data <=32'hFFB70018;
14'd6918:data <=32'hFFA00018;14'd6919:data <=32'hFF870022;14'd6920:data <=32'hFF74003D;
14'd6921:data <=32'hFF6B0061;14'd6922:data <=32'hFF700089;14'd6923:data <=32'hFF8400AD;
14'd6924:data <=32'hFFA200CC;14'd6925:data <=32'hFFC700E2;14'd6926:data <=32'hFFF000EE;
14'd6927:data <=32'h001B00F1;14'd6928:data <=32'h004500EB;14'd6929:data <=32'h006F00DB;
14'd6930:data <=32'h009500C3;14'd6931:data <=32'h00B500A1;14'd6932:data <=32'h00CD0076;
14'd6933:data <=32'h00D90048;14'd6934:data <=32'h00D50019;14'd6935:data <=32'h00C6FFEE;
14'd6936:data <=32'h00ACFFCD;14'd6937:data <=32'h008CFFB7;14'd6938:data <=32'h006BFFAC;
14'd6939:data <=32'h004FFFAC;14'd6940:data <=32'h0039FFB1;14'd6941:data <=32'h0026FFB9;
14'd6942:data <=32'h001AFFC2;14'd6943:data <=32'h000EFFCB;14'd6944:data <=32'h0005FFD5;
14'd6945:data <=32'hFFFCFFE1;14'd6946:data <=32'hFFF5FFEF;14'd6947:data <=32'hFFF40001;
14'd6948:data <=32'hFFF90014;14'd6949:data <=32'h00040026;14'd6950:data <=32'h00150034;
14'd6951:data <=32'h002B003D;14'd6952:data <=32'h0043003F;14'd6953:data <=32'h005D003B;
14'd6954:data <=32'h0075002F;14'd6955:data <=32'h008D001E;14'd6956:data <=32'h00A20007;
14'd6957:data <=32'h00B3FFEC;14'd6958:data <=32'h00BFFFC7;14'd6959:data <=32'h00C4FF9D;
14'd6960:data <=32'h00C0FF6F;14'd6961:data <=32'h00ACFF3F;14'd6962:data <=32'h008CFF10;
14'd6963:data <=32'h005CFEEC;14'd6964:data <=32'h0021FED4;14'd6965:data <=32'hFFE1FECF;
14'd6966:data <=32'hFFA3FEDC;14'd6967:data <=32'hFF6BFEF9;14'd6968:data <=32'hFF3FFF21;
14'd6969:data <=32'hFF22FF51;14'd6970:data <=32'hFF12FF82;14'd6971:data <=32'hFF0EFFB2;
14'd6972:data <=32'hFF15FFDD;14'd6973:data <=32'hFF210003;14'd6974:data <=32'hFF370023;
14'd6975:data <=32'hFF51003C;14'd6976:data <=32'hFF6AFFB1;14'd6977:data <=32'hFF4FFFC3;
14'd6978:data <=32'hFF35FFEB;14'd6979:data <=32'hFF47004C;14'd6980:data <=32'hFF820018;
14'd6981:data <=32'hFF840015;14'd6982:data <=32'hFF7F0015;14'd6983:data <=32'hFF76001A;
14'd6984:data <=32'hFF6C0029;14'd6985:data <=32'hFF68003F;14'd6986:data <=32'hFF6B0059;
14'd6987:data <=32'hFF770072;14'd6988:data <=32'hFF8A0087;14'd6989:data <=32'hFFA10095;
14'd6990:data <=32'hFFBA009C;14'd6991:data <=32'hFFD0009F;14'd6992:data <=32'hFFE4009F;
14'd6993:data <=32'hFFF8009D;14'd6994:data <=32'h000C0098;14'd6995:data <=32'h001E0091;
14'd6996:data <=32'h002F0086;14'd6997:data <=32'h003E0078;14'd6998:data <=32'h00470067;
14'd6999:data <=32'h004B0056;14'd7000:data <=32'h004A0049;14'd7001:data <=32'h00470040;
14'd7002:data <=32'h0043003B;14'd7003:data <=32'h00440039;14'd7004:data <=32'h00480037;
14'd7005:data <=32'h00510032;14'd7006:data <=32'h00590027;14'd7007:data <=32'h005E0018;
14'd7008:data <=32'h005C0005;14'd7009:data <=32'h0054FFF4;14'd7010:data <=32'h0044FFE7;
14'd7011:data <=32'h002FFFE0;14'd7012:data <=32'h001BFFE3;14'd7013:data <=32'h0009FFED;
14'd7014:data <=32'hFFFBFFFE;14'd7015:data <=32'hFFF60013;14'd7016:data <=32'hFFF80029;
14'd7017:data <=32'h0001003D;14'd7018:data <=32'h00110051;14'd7019:data <=32'h00270060;
14'd7020:data <=32'h0044006A;14'd7021:data <=32'h0066006D;14'd7022:data <=32'h008B0066;
14'd7023:data <=32'h00B20052;14'd7024:data <=32'h00D50032;14'd7025:data <=32'h00F00005;
14'd7026:data <=32'h00FCFFD0;14'd7027:data <=32'h00FAFF97;14'd7028:data <=32'h00E5FF61;
14'd7029:data <=32'h00C3FF32;14'd7030:data <=32'h0097FF10;14'd7031:data <=32'h0067FEFC;
14'd7032:data <=32'h0037FEF5;14'd7033:data <=32'h000AFEF6;14'd7034:data <=32'hFFE2FF00;
14'd7035:data <=32'hFFC1FF0E;14'd7036:data <=32'hFFA2FF1E;14'd7037:data <=32'hFF87FF32;
14'd7038:data <=32'hFF70FF49;14'd7039:data <=32'hFF60FF62;14'd7040:data <=32'hFF66FFA7;
14'd7041:data <=32'hFF5FFFBA;14'd7042:data <=32'hFF56FFBC;14'd7043:data <=32'hFF30FF6D;
14'd7044:data <=32'hFF49FF52;14'd7045:data <=32'hFF2EFF69;14'd7046:data <=32'hFF15FF88;
14'd7047:data <=32'hFEFFFFAC;14'd7048:data <=32'hFEF0FFD9;14'd7049:data <=32'hFEEC000D;
14'd7050:data <=32'hFEF70041;14'd7051:data <=32'hFF100072;14'd7052:data <=32'hFF370097;
14'd7053:data <=32'hFF6400AF;14'd7054:data <=32'hFF9200B9;14'd7055:data <=32'hFFBE00B5;
14'd7056:data <=32'hFFE100A7;14'd7057:data <=32'hFFFB0095;14'd7058:data <=32'h00100080;
14'd7059:data <=32'h001C0068;14'd7060:data <=32'h00210052;14'd7061:data <=32'h0021003D;
14'd7062:data <=32'h001A002A;14'd7063:data <=32'h000D001B;14'd7064:data <=32'hFFFD0014;
14'd7065:data <=32'hFFE90016;14'd7066:data <=32'hFFDA0021;14'd7067:data <=32'hFFD10035;
14'd7068:data <=32'hFFD20048;14'd7069:data <=32'hFFDD005C;14'd7070:data <=32'hFFF00069;
14'd7071:data <=32'h0006006E;14'd7072:data <=32'h001C0069;14'd7073:data <=32'h002D005D;
14'd7074:data <=32'h0037004D;14'd7075:data <=32'h003A003D;14'd7076:data <=32'h00360031;
14'd7077:data <=32'h00300028;14'd7078:data <=32'h00290025;14'd7079:data <=32'h00220025;
14'd7080:data <=32'h001D0028;14'd7081:data <=32'h001A002D;14'd7082:data <=32'h00190034;
14'd7083:data <=32'h001A003C;14'd7084:data <=32'h001F0046;14'd7085:data <=32'h00270051;
14'd7086:data <=32'h0036005A;14'd7087:data <=32'h004A005F;14'd7088:data <=32'h0062005F;
14'd7089:data <=32'h007B0057;14'd7090:data <=32'h00920046;14'd7091:data <=32'h00A2002F;
14'd7092:data <=32'h00AD0016;14'd7093:data <=32'h00AFFFFB;14'd7094:data <=32'h00ADFFE5;
14'd7095:data <=32'h00A8FFD3;14'd7096:data <=32'h00A3FFC4;14'd7097:data <=32'h00A3FFB5;
14'd7098:data <=32'h00A3FFA6;14'd7099:data <=32'h00A5FF90;14'd7100:data <=32'h00A1FF75;
14'd7101:data <=32'h0099FF57;14'd7102:data <=32'h0088FF38;14'd7103:data <=32'h006EFF1A;
14'd7104:data <=32'hFFBDFF2E;14'd7105:data <=32'hFFA7FF3A;14'd7106:data <=32'hFFADFF46;
14'd7107:data <=32'h002DFEFC;14'd7108:data <=32'h002DFEB6;14'd7109:data <=32'hFFEEFEA8;
14'd7110:data <=32'hFFAAFEA9;14'd7111:data <=32'hFF66FEBB;14'd7112:data <=32'hFF26FEDF;
14'd7113:data <=32'hFEEEFF16;14'd7114:data <=32'hFECAFF58;14'd7115:data <=32'hFEB9FFA2;
14'd7116:data <=32'hFEBEFFEC;14'd7117:data <=32'hFED6002C;14'd7118:data <=32'hFEFC005F;
14'd7119:data <=32'hFF290082;14'd7120:data <=32'hFF580097;14'd7121:data <=32'hFF8400A0;
14'd7122:data <=32'hFFAD009E;14'd7123:data <=32'hFFD20094;14'd7124:data <=32'hFFF20084;
14'd7125:data <=32'h0009006E;14'd7126:data <=32'h00170053;14'd7127:data <=32'h001E0037;
14'd7128:data <=32'h0019001D;14'd7129:data <=32'h000C0008;14'd7130:data <=32'hFFF9FFFC;
14'd7131:data <=32'hFFE6FFFA;14'd7132:data <=32'hFFD4FFFF;14'd7133:data <=32'hFFC9000B;
14'd7134:data <=32'hFFC30018;14'd7135:data <=32'hFFC40024;14'd7136:data <=32'hFFC7002C;
14'd7137:data <=32'hFFCA0031;14'd7138:data <=32'hFFCA0036;14'd7139:data <=32'hFFCA003B;
14'd7140:data <=32'hFFC80042;14'd7141:data <=32'hFFC8004E;14'd7142:data <=32'hFFCC005B;
14'd7143:data <=32'hFFD4006A;14'd7144:data <=32'hFFE10077;14'd7145:data <=32'hFFF30080;
14'd7146:data <=32'h00050084;14'd7147:data <=32'h00190084;14'd7148:data <=32'h002B0080;
14'd7149:data <=32'h003B007A;14'd7150:data <=32'h00490070;14'd7151:data <=32'h00560066;
14'd7152:data <=32'h00610059;14'd7153:data <=32'h0069004A;14'd7154:data <=32'h006D003A;
14'd7155:data <=32'h006D0029;14'd7156:data <=32'h0066001A;14'd7157:data <=32'h005B0012;
14'd7158:data <=32'h004E0011;14'd7159:data <=32'h00440019;14'd7160:data <=32'h00420028;
14'd7161:data <=32'h004A0039;14'd7162:data <=32'h005E0047;14'd7163:data <=32'h007D004E;
14'd7164:data <=32'h00A00048;14'd7165:data <=32'h00C40033;14'd7166:data <=32'h00E20012;
14'd7167:data <=32'h00F7FFE7;14'd7168:data <=32'h009AFF81;14'd7169:data <=32'h0097FF67;
14'd7170:data <=32'h0090FF69;14'd7171:data <=32'h00CBFFAC;14'd7172:data <=32'h00F2FF4E;
14'd7173:data <=32'h00D4FF1B;14'd7174:data <=32'h00A8FEEF;14'd7175:data <=32'h0072FECF;
14'd7176:data <=32'h0032FEBD;14'd7177:data <=32'hFFF0FEBE;14'd7178:data <=32'hFFB1FED1;
14'd7179:data <=32'hFF7EFEF3;14'd7180:data <=32'hFF58FF1E;14'd7181:data <=32'hFF3FFF4B;
14'd7182:data <=32'hFF36FF78;14'd7183:data <=32'hFF35FF9F;14'd7184:data <=32'hFF39FFC1;
14'd7185:data <=32'hFF40FFDF;14'd7186:data <=32'hFF4AFFF9;14'd7187:data <=32'hFF560011;
14'd7188:data <=32'hFF670027;14'd7189:data <=32'hFF7B0038;14'd7190:data <=32'hFF920043;
14'd7191:data <=32'hFFA80048;14'd7192:data <=32'hFFBD0046;14'd7193:data <=32'hFFCD0041;
14'd7194:data <=32'hFFD9003B;14'd7195:data <=32'hFFE20034;14'd7196:data <=32'hFFEA002D;
14'd7197:data <=32'hFFF00027;14'd7198:data <=32'hFFF8001D;14'd7199:data <=32'hFFFD0012;
14'd7200:data <=32'hFFFF0002;14'd7201:data <=32'hFFFAFFF1;14'd7202:data <=32'hFFEEFFE0;
14'd7203:data <=32'hFFD8FFD3;14'd7204:data <=32'hFFBEFFD0;14'd7205:data <=32'hFFA0FFD7;
14'd7206:data <=32'hFF85FFEA;14'd7207:data <=32'hFF720007;14'd7208:data <=32'hFF680028;
14'd7209:data <=32'hFF6A004C;14'd7210:data <=32'hFF75006D;14'd7211:data <=32'hFF88008B;
14'd7212:data <=32'hFFA300A2;14'd7213:data <=32'hFFC000B1;14'd7214:data <=32'hFFDF00BA;
14'd7215:data <=32'hFFFF00BB;14'd7216:data <=32'h001E00B7;14'd7217:data <=32'h003C00AB;
14'd7218:data <=32'h00540097;14'd7219:data <=32'h0065007E;14'd7220:data <=32'h006B0062;
14'd7221:data <=32'h00680049;14'd7222:data <=32'h005C0037;14'd7223:data <=32'h004D002F;
14'd7224:data <=32'h003E0031;14'd7225:data <=32'h0036003E;14'd7226:data <=32'h0036004F;
14'd7227:data <=32'h0043005F;14'd7228:data <=32'h005B006B;14'd7229:data <=32'h0077006D;
14'd7230:data <=32'h00960064;14'd7231:data <=32'h00B30052;14'd7232:data <=32'h0081006E;
14'd7233:data <=32'h00B00067;14'd7234:data <=32'h00C70051;14'd7235:data <=32'h00990013;
14'd7236:data <=32'h00CFFFCD;14'd7237:data <=32'h00C6FFB0;14'd7238:data <=32'h00B7FF94;
14'd7239:data <=32'h00A4FF79;14'd7240:data <=32'h008AFF65;14'd7241:data <=32'h006BFF59;
14'd7242:data <=32'h004CFF55;14'd7243:data <=32'h0033FF5A;14'd7244:data <=32'h0020FF64;
14'd7245:data <=32'h0015FF6D;14'd7246:data <=32'h000EFF72;14'd7247:data <=32'h000AFF72;
14'd7248:data <=32'h0002FF6C;14'd7249:data <=32'hFFF5FF64;14'd7250:data <=32'hFFE1FF5F;
14'd7251:data <=32'hFFC9FF60;14'd7252:data <=32'hFFB0FF68;14'd7253:data <=32'hFF97FF76;
14'd7254:data <=32'hFF84FF8A;14'd7255:data <=32'hFF77FFA3;14'd7256:data <=32'hFF6FFFBD;
14'd7257:data <=32'hFF6CFFD7;14'd7258:data <=32'hFF6EFFF1;14'd7259:data <=32'hFF76000B;
14'd7260:data <=32'hFF840023;14'd7261:data <=32'hFF990039;14'd7262:data <=32'hFFB40046;
14'd7263:data <=32'hFFD30049;14'd7264:data <=32'hFFF20041;14'd7265:data <=32'h000C002F;
14'd7266:data <=32'h001D0012;14'd7267:data <=32'h0021FFF1;14'd7268:data <=32'h0018FFD1;
14'd7269:data <=32'h0003FFB8;14'd7270:data <=32'hFFE5FFA8;14'd7271:data <=32'hFFC4FFA3;
14'd7272:data <=32'hFFA5FFAA;14'd7273:data <=32'hFF8AFFB9;14'd7274:data <=32'hFF74FFCE;
14'd7275:data <=32'hFF64FFE7;14'd7276:data <=32'hFF5B0002;14'd7277:data <=32'hFF57001E;
14'd7278:data <=32'hFF57003A;14'd7279:data <=32'hFF5E0057;14'd7280:data <=32'hFF6A0073;
14'd7281:data <=32'hFF7C008B;14'd7282:data <=32'hFF93009E;14'd7283:data <=32'hFFAB00AA;
14'd7284:data <=32'hFFC300B1;14'd7285:data <=32'hFFD900B2;14'd7286:data <=32'hFFEB00B2;
14'd7287:data <=32'hFFF900B3;14'd7288:data <=32'h000700B7;14'd7289:data <=32'h001800BD;
14'd7290:data <=32'h002E00C4;14'd7291:data <=32'h004B00C8;14'd7292:data <=32'h006C00C5;
14'd7293:data <=32'h009100B7;14'd7294:data <=32'h00B1009F;14'd7295:data <=32'h00CA0080;
14'd7296:data <=32'hFFE40083;14'd7297:data <=32'h000800AE;14'd7298:data <=32'h004300BC;
14'd7299:data <=32'h00C30039;14'd7300:data <=32'h00EDFFE9;14'd7301:data <=32'h00D6FFC6;
14'd7302:data <=32'h00BBFFAB;14'd7303:data <=32'h009CFF98;14'd7304:data <=32'h007BFF8E;
14'd7305:data <=32'h0059FF8C;14'd7306:data <=32'h003DFF97;14'd7307:data <=32'h0027FFAB;
14'd7308:data <=32'h001EFFC1;14'd7309:data <=32'h0023FFD9;14'd7310:data <=32'h0031FFE7;
14'd7311:data <=32'h0047FFEA;14'd7312:data <=32'h005BFFE1;14'd7313:data <=32'h006AFFCD;
14'd7314:data <=32'h0070FFB1;14'd7315:data <=32'h0069FF96;14'd7316:data <=32'h005AFF7B;
14'd7317:data <=32'h0043FF68;14'd7318:data <=32'h0028FF5D;14'd7319:data <=32'h000CFF57;
14'd7320:data <=32'hFFEFFF58;14'd7321:data <=32'hFFD3FF5F;14'd7322:data <=32'hFFB9FF6C;
14'd7323:data <=32'hFFA1FF80;14'd7324:data <=32'hFF8FFF99;14'd7325:data <=32'hFF85FFB8;
14'd7326:data <=32'hFF85FFD7;14'd7327:data <=32'hFF90FFF3;14'd7328:data <=32'hFFA4000B;
14'd7329:data <=32'hFFBC0017;14'd7330:data <=32'hFFD5001A;14'd7331:data <=32'hFFEA0012;
14'd7332:data <=32'hFFF90005;14'd7333:data <=32'h0000FFF5;14'd7334:data <=32'h0000FFE6;
14'd7335:data <=32'hFFFDFFD8;14'd7336:data <=32'hFFF7FFCE;14'd7337:data <=32'hFFEFFFC6;
14'd7338:data <=32'hFFE7FFC0;14'd7339:data <=32'hFFDFFFB8;14'd7340:data <=32'hFFD4FFAF;
14'd7341:data <=32'hFFC5FFA8;14'd7342:data <=32'hFFB1FFA3;14'd7343:data <=32'hFF99FFA3;
14'd7344:data <=32'hFF7FFFA9;14'd7345:data <=32'hFF65FFB7;14'd7346:data <=32'hFF4DFFCA;
14'd7347:data <=32'hFF38FFE3;14'd7348:data <=32'hFF270002;14'd7349:data <=32'hFF1C0023;
14'd7350:data <=32'hFF150049;14'd7351:data <=32'hFF140075;14'd7352:data <=32'hFF1B00A4;
14'd7353:data <=32'hFF2D00D5;14'd7354:data <=32'hFF4F0106;14'd7355:data <=32'hFF7E0131;
14'd7356:data <=32'hFFBC0150;14'd7357:data <=32'h0002015C;14'd7358:data <=32'h00490156;
14'd7359:data <=32'h008D013B;14'd7360:data <=32'hFFDD006B;14'd7361:data <=32'hFFE50091;
14'd7362:data <=32'h000300C4;14'd7363:data <=32'h00A300FD;14'd7364:data <=32'h00F400A4;
14'd7365:data <=32'h00FB006F;14'd7366:data <=32'h00F9003C;14'd7367:data <=32'h00EA000F;
14'd7368:data <=32'h00D3FFE9;14'd7369:data <=32'h00B4FFCC;14'd7370:data <=32'h0092FFBB;
14'd7371:data <=32'h0070FFB8;14'd7372:data <=32'h0054FFC0;14'd7373:data <=32'h0042FFD0;
14'd7374:data <=32'h003DFFE0;14'd7375:data <=32'h0041FFEE;14'd7376:data <=32'h004CFFF4;
14'd7377:data <=32'h0058FFF1;14'd7378:data <=32'h0060FFE6;14'd7379:data <=32'h0064FFD8;
14'd7380:data <=32'h0061FFC9;14'd7381:data <=32'h005AFFBD;14'd7382:data <=32'h0051FFB3;
14'd7383:data <=32'h0047FFAD;14'd7384:data <=32'h003EFFA8;14'd7385:data <=32'h0035FFA2;
14'd7386:data <=32'h002CFF9D;14'd7387:data <=32'h001FFF9A;14'd7388:data <=32'h0011FF99;
14'd7389:data <=32'h0005FF9C;14'd7390:data <=32'hFFFAFFA2;14'd7391:data <=32'hFFF2FFAB;
14'd7392:data <=32'hFFEEFFB2;14'd7393:data <=32'hFFEDFFBA;14'd7394:data <=32'hFFEEFFBD;
14'd7395:data <=32'hFFEEFFBD;14'd7396:data <=32'hFFEAFFBC;14'd7397:data <=32'hFFE4FFBD;
14'd7398:data <=32'hFFDCFFC0;14'd7399:data <=32'hFFD6FFC7;14'd7400:data <=32'hFFD2FFD3;
14'd7401:data <=32'hFFD6FFE0;14'd7402:data <=32'hFFDFFFEA;14'd7403:data <=32'hFFEEFFED;
14'd7404:data <=32'h0000FFE9;14'd7405:data <=32'h000DFFDC;14'd7406:data <=32'h0016FFC7;
14'd7407:data <=32'h0016FFAD;14'd7408:data <=32'h000CFF93;14'd7409:data <=32'hFFF9FF7B;
14'd7410:data <=32'hFFDDFF68;14'd7411:data <=32'hFFBBFF5A;14'd7412:data <=32'hFF93FF55;
14'd7413:data <=32'hFF67FF5A;14'd7414:data <=32'hFF3AFF6A;14'd7415:data <=32'hFF0EFF86;
14'd7416:data <=32'hFEE5FFB0;14'd7417:data <=32'hFEC5FFE7;14'd7418:data <=32'hFEB5002B;
14'd7419:data <=32'hFEB70073;14'd7420:data <=32'hFECE00BB;14'd7421:data <=32'hFEF800FA;
14'd7422:data <=32'hFF34012A;14'd7423:data <=32'hFF760147;14'd7424:data <=32'hFF8300BA;
14'd7425:data <=32'hFF9400E0;14'd7426:data <=32'hFF9C0103;14'd7427:data <=32'hFF93012D;
14'd7428:data <=32'hFFF80107;14'd7429:data <=32'h001B00FD;14'd7430:data <=32'h003C00EE;
14'd7431:data <=32'h005900DC;14'd7432:data <=32'h007200C5;14'd7433:data <=32'h008400AC;
14'd7434:data <=32'h00900092;14'd7435:data <=32'h0096007A;14'd7436:data <=32'h00990067;
14'd7437:data <=32'h009E0056;14'd7438:data <=32'h00A30047;14'd7439:data <=32'h00AA0034;
14'd7440:data <=32'h00B1001D;14'd7441:data <=32'h00B40002;14'd7442:data <=32'h00AEFFE4;
14'd7443:data <=32'h009FFFC7;14'd7444:data <=32'h0087FFB0;14'd7445:data <=32'h006AFFA1;
14'd7446:data <=32'h004CFF9E;14'd7447:data <=32'h0031FFA3;14'd7448:data <=32'h001EFFB0;
14'd7449:data <=32'h0010FFC0;14'd7450:data <=32'h000AFFD1;14'd7451:data <=32'h000AFFDF;
14'd7452:data <=32'h000DFFEC;14'd7453:data <=32'h0014FFF5;14'd7454:data <=32'h001EFFFC;
14'd7455:data <=32'h002A0000;14'd7456:data <=32'h0039FFFE;14'd7457:data <=32'h0046FFF8;
14'd7458:data <=32'h0051FFE9;14'd7459:data <=32'h0059FFD6;14'd7460:data <=32'h0057FFC1;
14'd7461:data <=32'h004EFFAC;14'd7462:data <=32'h003DFF9A;14'd7463:data <=32'h0027FF92;
14'd7464:data <=32'h0011FF92;14'd7465:data <=32'hFFFEFF9C;14'd7466:data <=32'hFFF3FFA9;
14'd7467:data <=32'hFFF0FFB7;14'd7468:data <=32'hFFF5FFC4;14'd7469:data <=32'hFFFFFFC9;
14'd7470:data <=32'h000BFFC7;14'd7471:data <=32'h0014FFBE;14'd7472:data <=32'h0018FFB0;
14'd7473:data <=32'h0018FF9F;14'd7474:data <=32'h0010FF8E;14'd7475:data <=32'h0004FF7D;
14'd7476:data <=32'hFFF3FF6D;14'd7477:data <=32'hFFDDFF5E;14'd7478:data <=32'hFFC0FF54;
14'd7479:data <=32'hFF9FFF51;14'd7480:data <=32'hFF78FF56;14'd7481:data <=32'hFF52FF66;
14'd7482:data <=32'hFF2DFF82;14'd7483:data <=32'hFF11FFA9;14'd7484:data <=32'hFEFFFFD6;
14'd7485:data <=32'hFEFC0005;14'd7486:data <=32'hFF060032;14'd7487:data <=32'hFF170057;
14'd7488:data <=32'hFECA003A;14'd7489:data <=32'hFEC4007D;14'd7490:data <=32'hFED500A6;
14'd7491:data <=32'hFF1B004C;14'd7492:data <=32'hFF53003E;14'd7493:data <=32'hFF4F0052;
14'd7494:data <=32'hFF4F006C;14'd7495:data <=32'hFF55008B;14'd7496:data <=32'hFF6300A9;
14'd7497:data <=32'hFF7900C5;14'd7498:data <=32'hFF9400DD;14'd7499:data <=32'hFFB500F2;
14'd7500:data <=32'hFFDA0101;14'd7501:data <=32'h0003010B;14'd7502:data <=32'h0033010E;
14'd7503:data <=32'h00660104;14'd7504:data <=32'h009800EC;14'd7505:data <=32'h00C300C7;
14'd7506:data <=32'h00E30094;14'd7507:data <=32'h00F4005A;14'd7508:data <=32'h00F20020;
14'd7509:data <=32'h00DEFFEC;14'd7510:data <=32'h00BEFFC2;14'd7511:data <=32'h0097FFA8;
14'd7512:data <=32'h006EFF9A;14'd7513:data <=32'h0049FF99;14'd7514:data <=32'h0029FFA1;
14'd7515:data <=32'h000EFFB0;14'd7516:data <=32'hFFFAFFC3;14'd7517:data <=32'hFFECFFDA;
14'd7518:data <=32'hFFE6FFF3;14'd7519:data <=32'hFFEA000D;14'd7520:data <=32'hFFF40024;
14'd7521:data <=32'h00070036;14'd7522:data <=32'h001F003F;14'd7523:data <=32'h00380040;
14'd7524:data <=32'h00510038;14'd7525:data <=32'h00630029;14'd7526:data <=32'h00710015;
14'd7527:data <=32'h00750000;14'd7528:data <=32'h0075FFEF;14'd7529:data <=32'h0073FFE0;
14'd7530:data <=32'h0070FFD6;14'd7531:data <=32'h006EFFCC;14'd7532:data <=32'h0070FFC1;
14'd7533:data <=32'h0070FFB2;14'd7534:data <=32'h0071FF9F;14'd7535:data <=32'h006AFF8B;
14'd7536:data <=32'h005FFF75;14'd7537:data <=32'h004CFF61;14'd7538:data <=32'h0034FF50;
14'd7539:data <=32'h0019FF48;14'd7540:data <=32'hFFFDFF44;14'd7541:data <=32'hFFE2FF46;
14'd7542:data <=32'hFFC9FF4C;14'd7543:data <=32'hFFB1FF55;14'd7544:data <=32'hFF9BFF62;
14'd7545:data <=32'hFF86FF73;14'd7546:data <=32'hFF75FF89;14'd7547:data <=32'hFF69FFA2;
14'd7548:data <=32'hFF65FFBD;14'd7549:data <=32'hFF6BFFD7;14'd7550:data <=32'hFF76FFE9;
14'd7551:data <=32'hFF85FFF3;14'd7552:data <=32'hFF1BFF52;14'd7553:data <=32'hFEE8FF77;
14'd7554:data <=32'hFEDAFFAE;14'd7555:data <=32'hFF7AFFDE;14'd7556:data <=32'hFFA8FFB4;
14'd7557:data <=32'hFF8DFFAE;14'd7558:data <=32'hFF6FFFB3;14'd7559:data <=32'hFF50FFC3;
14'd7560:data <=32'hFF37FFDE;14'd7561:data <=32'hFF240000;14'd7562:data <=32'hFF1A0026;
14'd7563:data <=32'hFF170051;14'd7564:data <=32'hFF1E007E;14'd7565:data <=32'hFF3000AC;
14'd7566:data <=32'hFF4F00D8;14'd7567:data <=32'hFF7B00FC;14'd7568:data <=32'hFFB20113;
14'd7569:data <=32'hFFEE0119;14'd7570:data <=32'h0029010F;14'd7571:data <=32'h005C00F5;
14'd7572:data <=32'h008500CE;14'd7573:data <=32'h009D00A2;14'd7574:data <=32'h00A70074;
14'd7575:data <=32'h00A6004C;14'd7576:data <=32'h009C0029;14'd7577:data <=32'h008E000E;
14'd7578:data <=32'h007DFFF8;14'd7579:data <=32'h006BFFE7;14'd7580:data <=32'h0055FFDA;
14'd7581:data <=32'h0040FFD3;14'd7582:data <=32'h0028FFD2;14'd7583:data <=32'h0011FFD8;
14'd7584:data <=32'hFFFFFFE3;14'd7585:data <=32'hFFF2FFF5;14'd7586:data <=32'hFFEB0008;
14'd7587:data <=32'hFFEB001C;14'd7588:data <=32'hFFF0002E;14'd7589:data <=32'hFFF9003D;
14'd7590:data <=32'h0004004A;14'd7591:data <=32'h00120055;14'd7592:data <=32'h0022005F;
14'd7593:data <=32'h00350068;14'd7594:data <=32'h004D006F;14'd7595:data <=32'h006B0070;
14'd7596:data <=32'h008E0069;14'd7597:data <=32'h00B10057;14'd7598:data <=32'h00D40039;
14'd7599:data <=32'h00EC000E;14'd7600:data <=32'h00F8FFDD;14'd7601:data <=32'h00F6FFA7;
14'd7602:data <=32'h00E5FF74;14'd7603:data <=32'h00C7FF46;14'd7604:data <=32'h00A0FF23;
14'd7605:data <=32'h0073FF0B;14'd7606:data <=32'h0044FEFE;14'd7607:data <=32'h0014FEFB;
14'd7608:data <=32'hFFE6FF03;14'd7609:data <=32'hFFBCFF14;14'd7610:data <=32'hFF97FF2E;
14'd7611:data <=32'hFF7CFF51;14'd7612:data <=32'hFF6CFF78;14'd7613:data <=32'hFF6AFFA0;
14'd7614:data <=32'hFF74FFC3;14'd7615:data <=32'hFF88FFDC;14'd7616:data <=32'hFFCFFF5F;
14'd7617:data <=32'hFFB3FF53;14'd7618:data <=32'hFF89FF60;14'd7619:data <=32'hFF78FFC2;
14'd7620:data <=32'hFFB4FFA2;14'd7621:data <=32'hFFA7FF9C;14'd7622:data <=32'hFF96FF9B;
14'd7623:data <=32'hFF80FFA1;14'd7624:data <=32'hFF6EFFAF;14'd7625:data <=32'hFF5FFFC0;
14'd7626:data <=32'hFF53FFD4;14'd7627:data <=32'hFF4AFFE9;14'd7628:data <=32'hFF430002;
14'd7629:data <=32'hFF40001E;14'd7630:data <=32'hFF43003D;14'd7631:data <=32'hFF50005C;
14'd7632:data <=32'hFF640078;14'd7633:data <=32'hFF7F008D;14'd7634:data <=32'hFF9D0099;
14'd7635:data <=32'hFFBE009C;14'd7636:data <=32'hFFD80096;14'd7637:data <=32'hFFEB008B;
14'd7638:data <=32'hFFF90081;14'd7639:data <=32'h00000078;14'd7640:data <=32'h00070072;
14'd7641:data <=32'h000F0070;14'd7642:data <=32'h0019006D;14'd7643:data <=32'h00260068;
14'd7644:data <=32'h0033005E;14'd7645:data <=32'h003E0050;14'd7646:data <=32'h00450040;
14'd7647:data <=32'h0046002D;14'd7648:data <=32'h0041001C;14'd7649:data <=32'h0038000D;
14'd7650:data <=32'h002C0004;14'd7651:data <=32'h001EFFFD;14'd7652:data <=32'h000EFFFB;
14'd7653:data <=32'hFFFEFFFD;14'd7654:data <=32'hFFED0004;14'd7655:data <=32'hFFDE0011;
14'd7656:data <=32'hFFD00026;14'd7657:data <=32'hFFC90041;14'd7658:data <=32'hFFCC0062;
14'd7659:data <=32'hFFDA0085;14'd7660:data <=32'hFFF700A4;14'd7661:data <=32'h002000BB;
14'd7662:data <=32'h005200C3;14'd7663:data <=32'h008600BC;14'd7664:data <=32'h00B700A5;
14'd7665:data <=32'h00E00081;14'd7666:data <=32'h00FC0053;14'd7667:data <=32'h010C0021;
14'd7668:data <=32'h0110FFEE;14'd7669:data <=32'h0108FFBD;14'd7670:data <=32'h00F7FF92;
14'd7671:data <=32'h00DFFF6B;14'd7672:data <=32'h00C1FF4A;14'd7673:data <=32'h009CFF30;
14'd7674:data <=32'h0075FF1F;14'd7675:data <=32'h004BFF19;14'd7676:data <=32'h0023FF1D;
14'd7677:data <=32'h0003FF29;14'd7678:data <=32'hFFEBFF3B;14'd7679:data <=32'hFFDBFF4C;
14'd7680:data <=32'hFFD5FF92;14'd7681:data <=32'hFFDBFF93;14'd7682:data <=32'hFFD6FF80;
14'd7683:data <=32'hFFBDFF24;14'd7684:data <=32'hFFDBFF09;14'd7685:data <=32'hFFB2FF0D;
14'd7686:data <=32'hFF88FF1B;14'd7687:data <=32'hFF61FF35;14'd7688:data <=32'hFF42FF59;
14'd7689:data <=32'hFF2FFF82;14'd7690:data <=32'hFF28FFAC;14'd7691:data <=32'hFF29FFD2;
14'd7692:data <=32'hFF32FFF7;14'd7693:data <=32'hFF400014;14'd7694:data <=32'hFF530030;
14'd7695:data <=32'hFF690044;14'd7696:data <=32'hFF840053;14'd7697:data <=32'hFFA0005A;
14'd7698:data <=32'hFFBD0058;14'd7699:data <=32'hFFD5004C;14'd7700:data <=32'hFFE4003A;
14'd7701:data <=32'hFFE70024;14'd7702:data <=32'hFFE20012;14'd7703:data <=32'hFFD40008;
14'd7704:data <=32'hFFC10007;14'd7705:data <=32'hFFB20010;14'd7706:data <=32'hFFA80020;
14'd7707:data <=32'hFFA70035;14'd7708:data <=32'hFFAE0047;14'd7709:data <=32'hFFBB0057;
14'd7710:data <=32'hFFCC005F;14'd7711:data <=32'hFFDD0063;14'd7712:data <=32'hFFEE0062;
14'd7713:data <=32'hFFFB005C;14'd7714:data <=32'h00070054;14'd7715:data <=32'h000F004B;
14'd7716:data <=32'h0016003E;14'd7717:data <=32'h00160031;14'd7718:data <=32'h00120024;
14'd7719:data <=32'h0008001A;14'd7720:data <=32'hFFF90016;14'd7721:data <=32'hFFE70019;
14'd7722:data <=32'hFFD60024;14'd7723:data <=32'hFFCB0039;14'd7724:data <=32'hFFC70052;
14'd7725:data <=32'hFFCE006D;14'd7726:data <=32'hFFE10085;14'd7727:data <=32'hFFF90097;
14'd7728:data <=32'h001600A1;14'd7729:data <=32'h003400A0;14'd7730:data <=32'h004F009B;
14'd7731:data <=32'h00660091;14'd7732:data <=32'h007A0084;14'd7733:data <=32'h008A0078;
14'd7734:data <=32'h009C006B;14'd7735:data <=32'h00AE005D;14'd7736:data <=32'h00BF0048;
14'd7737:data <=32'h00CF0032;14'd7738:data <=32'h00DB0017;14'd7739:data <=32'h00E3FFF9;
14'd7740:data <=32'h00E5FFDA;14'd7741:data <=32'h00E4FFBC;14'd7742:data <=32'h00E0FF9E;
14'd7743:data <=32'h00DBFF80;14'd7744:data <=32'h0024FF60;14'd7745:data <=32'h0020FF67;
14'd7746:data <=32'h0033FF6C;14'd7747:data <=32'h00C8FF37;14'd7748:data <=32'h00E2FEEC;
14'd7749:data <=32'h00A7FEBF;14'd7750:data <=32'h0062FEA3;14'd7751:data <=32'h0016FE99;
14'd7752:data <=32'hFFCCFEA5;14'd7753:data <=32'hFF8BFEC4;14'd7754:data <=32'hFF58FEEF;
14'd7755:data <=32'hFF33FF21;14'd7756:data <=32'hFF1CFF58;14'd7757:data <=32'hFF13FF8F;
14'd7758:data <=32'hFF14FFC2;14'd7759:data <=32'hFF22FFF2;14'd7760:data <=32'hFF3A001C;
14'd7761:data <=32'hFF5B003D;14'd7762:data <=32'hFF82004F;14'd7763:data <=32'hFFAA0055;
14'd7764:data <=32'hFFCE004D;14'd7765:data <=32'hFFE9003A;14'd7766:data <=32'hFFF80020;
14'd7767:data <=32'hFFFA0007;14'd7768:data <=32'hFFF3FFF4;14'd7769:data <=32'hFFE4FFE7;
14'd7770:data <=32'hFFD6FFE2;14'd7771:data <=32'hFFC8FFE6;14'd7772:data <=32'hFFBEFFEC;
14'd7773:data <=32'hFFB9FFF4;14'd7774:data <=32'hFFB4FFFB;14'd7775:data <=32'hFFB20002;
14'd7776:data <=32'hFFB00007;14'd7777:data <=32'hFFAD000F;14'd7778:data <=32'hFFAB0017;
14'd7779:data <=32'hFFAB0022;14'd7780:data <=32'hFFAC002C;14'd7781:data <=32'hFFB00034;
14'd7782:data <=32'hFFB6003C;14'd7783:data <=32'hFFBC0041;14'd7784:data <=32'hFFC10045;
14'd7785:data <=32'hFFC4004B;14'd7786:data <=32'hFFC60051;14'd7787:data <=32'hFFCA0059;
14'd7788:data <=32'hFFD10063;14'd7789:data <=32'hFFDC006C;14'd7790:data <=32'hFFEA0073;
14'd7791:data <=32'hFFFB0073;14'd7792:data <=32'h000B006E;14'd7793:data <=32'h00160065;
14'd7794:data <=32'h001B0059;14'd7795:data <=32'h0018004F;14'd7796:data <=32'h0010004B;
14'd7797:data <=32'h0006004F;14'd7798:data <=32'hFFFF005B;14'd7799:data <=32'hFFFE006E;
14'd7800:data <=32'h00070084;14'd7801:data <=32'h00190098;14'd7802:data <=32'h003200A8;
14'd7803:data <=32'h005300B3;14'd7804:data <=32'h007800B5;14'd7805:data <=32'h00A000B1;
14'd7806:data <=32'h00CB00A2;14'd7807:data <=32'h00F50089;14'd7808:data <=32'h00B0FFF4;
14'd7809:data <=32'h00C2FFE9;14'd7810:data <=32'h00CCFFED;14'd7811:data <=32'h010A003D;
14'd7812:data <=32'h015AFFE7;14'd7813:data <=32'h0151FFA0;14'd7814:data <=32'h0135FF5D;
14'd7815:data <=32'h0108FF25;14'd7816:data <=32'h00D2FEFD;14'd7817:data <=32'h0096FEE7;
14'd7818:data <=32'h005DFEDF;14'd7819:data <=32'h0028FEE2;14'd7820:data <=32'hFFF8FEEF;
14'd7821:data <=32'hFFCEFF02;14'd7822:data <=32'hFFAAFF1C;14'd7823:data <=32'hFF8CFF3C;
14'd7824:data <=32'hFF78FF60;14'd7825:data <=32'hFF6DFF85;14'd7826:data <=32'hFF6CFFA9;
14'd7827:data <=32'hFF76FFC7;14'd7828:data <=32'hFF84FFDF;14'd7829:data <=32'hFF94FFEE;
14'd7830:data <=32'hFFA3FFF6;14'd7831:data <=32'hFFAFFFFA;14'd7832:data <=32'hFFB5FFFC;
14'd7833:data <=32'hFFBB0000;14'd7834:data <=32'hFFC10005;14'd7835:data <=32'hFFCA000C;
14'd7836:data <=32'hFFD7000F;14'd7837:data <=32'hFFE5000D;14'd7838:data <=32'hFFF20006;
14'd7839:data <=32'hFFFBFFF8;14'd7840:data <=32'hFFFEFFE6;14'd7841:data <=32'hFFF9FFD3;
14'd7842:data <=32'hFFEDFFC3;14'd7843:data <=32'hFFDAFFB8;14'd7844:data <=32'hFFC5FFB4;
14'd7845:data <=32'hFFAEFFB7;14'd7846:data <=32'hFF99FFBF;14'd7847:data <=32'hFF85FFCE;
14'd7848:data <=32'hFF75FFE0;14'd7849:data <=32'hFF68FFF6;14'd7850:data <=32'hFF60000F;
14'd7851:data <=32'hFF5F002D;14'd7852:data <=32'hFF66004C;14'd7853:data <=32'hFF740069;
14'd7854:data <=32'hFF8C0082;14'd7855:data <=32'hFFAA0091;14'd7856:data <=32'hFFCA0095;
14'd7857:data <=32'hFFE8008E;14'd7858:data <=32'hFFFE007E;14'd7859:data <=32'h00090069;
14'd7860:data <=32'h00090055;14'd7861:data <=32'h00010046;14'd7862:data <=32'hFFF30042;
14'd7863:data <=32'hFFE50047;14'd7864:data <=32'hFFDA0054;14'd7865:data <=32'hFFD50068;
14'd7866:data <=32'hFFD7007E;14'd7867:data <=32'hFFE20094;14'd7868:data <=32'hFFF400AA;
14'd7869:data <=32'h000C00BD;14'd7870:data <=32'h002B00CD;14'd7871:data <=32'h005200D6;
14'd7872:data <=32'h002C00C0;14'd7873:data <=32'h005F00DA;14'd7874:data <=32'h008500DB;
14'd7875:data <=32'h007800A4;14'd7876:data <=32'h00D60073;14'd7877:data <=32'h00E4004C;
14'd7878:data <=32'h00E70023;14'd7879:data <=32'h00E0FFFB;14'd7880:data <=32'h00D1FFDE;
14'd7881:data <=32'h00BFFFC8;14'd7882:data <=32'h00B0FFB9;14'd7883:data <=32'h00A3FFAD;
14'd7884:data <=32'h0098FFA1;14'd7885:data <=32'h008FFF94;14'd7886:data <=32'h0083FF85;
14'd7887:data <=32'h0075FF75;14'd7888:data <=32'h0061FF68;14'd7889:data <=32'h004CFF5E;
14'd7890:data <=32'h0036FF5A;14'd7891:data <=32'h0021FF57;14'd7892:data <=32'h000CFF58;
14'd7893:data <=32'hFFF5FF57;14'd7894:data <=32'hFFDFFF5B;14'd7895:data <=32'hFFC5FF63;
14'd7896:data <=32'hFFACFF72;14'd7897:data <=32'hFF96FF89;14'd7898:data <=32'hFF85FFA9;
14'd7899:data <=32'hFF80FFCB;14'd7900:data <=32'hFF86FFEE;14'd7901:data <=32'hFF9A000C;
14'd7902:data <=32'hFFB60021;14'd7903:data <=32'hFFD5002A;14'd7904:data <=32'hFFF50025;
14'd7905:data <=32'h000F0016;14'd7906:data <=32'h00210001;14'd7907:data <=32'h0029FFE5;
14'd7908:data <=32'h0029FFCC;14'd7909:data <=32'h001FFFB3;14'd7910:data <=32'h000FFF9E;
14'd7911:data <=32'hFFFBFF8D;14'd7912:data <=32'hFFE0FF82;14'd7913:data <=32'hFFC3FF7D;
14'd7914:data <=32'hFFA3FF81;14'd7915:data <=32'hFF85FF8D;14'd7916:data <=32'hFF6AFFA2;
14'd7917:data <=32'hFF55FFBE;14'd7918:data <=32'hFF4AFFDF;14'd7919:data <=32'hFF490000;
14'd7920:data <=32'hFF50001C;14'd7921:data <=32'hFF5D0033;14'd7922:data <=32'hFF6C0041;
14'd7923:data <=32'hFF77004B;14'd7924:data <=32'hFF7F0052;14'd7925:data <=32'hFF840059;
14'd7926:data <=32'hFF850065;14'd7927:data <=32'hFF880074;14'd7928:data <=32'hFF8F0086;
14'd7929:data <=32'hFF9A009C;14'd7930:data <=32'hFFAD00AE;14'd7931:data <=32'hFFC300BD;
14'd7932:data <=32'hFFDE00C7;14'd7933:data <=32'hFFF800CC;14'd7934:data <=32'h001400CE;
14'd7935:data <=32'h002F00CB;14'd7936:data <=32'hFF6D007E;14'd7937:data <=32'hFF7C00C6;
14'd7938:data <=32'hFFB100F5;14'd7939:data <=32'h005800A8;14'd7940:data <=32'h00AB0078;
14'd7941:data <=32'h00AC0051;14'd7942:data <=32'h00A3002E;14'd7943:data <=32'h00910011;
14'd7944:data <=32'h00780002;14'd7945:data <=32'h00600000;14'd7946:data <=32'h004D0008;
14'd7947:data <=32'h00450016;14'd7948:data <=32'h00490025;14'd7949:data <=32'h0056002F;
14'd7950:data <=32'h00680032;14'd7951:data <=32'h007B002C;14'd7952:data <=32'h008D001E;
14'd7953:data <=32'h009B000B;14'd7954:data <=32'h00A6FFF4;14'd7955:data <=32'h00AAFFD9;
14'd7956:data <=32'h00AAFFBC;14'd7957:data <=32'h00A2FF9C;14'd7958:data <=32'h0091FF7E;
14'd7959:data <=32'h0077FF61;14'd7960:data <=32'h0054FF4C;14'd7961:data <=32'h002AFF42;
14'd7962:data <=32'h0001FF48;14'd7963:data <=32'hFFDBFF58;14'd7964:data <=32'hFFBDFF75;
14'd7965:data <=32'hFFACFF96;14'd7966:data <=32'hFFA8FFB9;14'd7967:data <=32'hFFAFFFD7;
14'd7968:data <=32'hFFBDFFEE;14'd7969:data <=32'hFFD0FFFC;14'd7970:data <=32'hFFE40003;
14'd7971:data <=32'hFFF50004;14'd7972:data <=32'h00050001;14'd7973:data <=32'h0013FFFB;
14'd7974:data <=32'h001EFFF1;14'd7975:data <=32'h0028FFE3;14'd7976:data <=32'h002FFFD1;
14'd7977:data <=32'h0030FFBE;14'd7978:data <=32'h002CFFA9;14'd7979:data <=32'h0021FF94;
14'd7980:data <=32'h0011FF83;14'd7981:data <=32'hFFFCFF75;14'd7982:data <=32'hFFE6FF6D;
14'd7983:data <=32'hFFCEFF6A;14'd7984:data <=32'hFFB7FF6A;14'd7985:data <=32'hFFA0FF6B;
14'd7986:data <=32'hFF87FF6D;14'd7987:data <=32'hFF6AFF72;14'd7988:data <=32'hFF4AFF7F;
14'd7989:data <=32'hFF28FF92;14'd7990:data <=32'hFF06FFB2;14'd7991:data <=32'hFEEAFFDE;
14'd7992:data <=32'hFEDA0012;14'd7993:data <=32'hFED7004E;14'd7994:data <=32'hFEE6008A;
14'd7995:data <=32'hFF0300C0;14'd7996:data <=32'hFF2D00EC;14'd7997:data <=32'hFF5F010C;
14'd7998:data <=32'hFF940120;14'd7999:data <=32'hFFCB0128;14'd8000:data <=32'hFF760025;
14'd8001:data <=32'hFF5E0059;14'd8002:data <=32'hFF6300A2;14'd8003:data <=32'hFFF7011C;
14'd8004:data <=32'h006900F1;14'd8005:data <=32'h008800C4;14'd8006:data <=32'h00980095;
14'd8007:data <=32'h00980067;14'd8008:data <=32'h00890040;14'd8009:data <=32'h00720029;
14'd8010:data <=32'h0059001E;14'd8011:data <=32'h0044001F;14'd8012:data <=32'h00370028;
14'd8013:data <=32'h00340034;14'd8014:data <=32'h0038003D;14'd8015:data <=32'h00410043;
14'd8016:data <=32'h004D0045;14'd8017:data <=32'h00590042;14'd8018:data <=32'h0065003E;
14'd8019:data <=32'h00710036;14'd8020:data <=32'h007E002A;14'd8021:data <=32'h0089001A;
14'd8022:data <=32'h00920005;14'd8023:data <=32'h0093FFEB;14'd8024:data <=32'h008EFFD3;
14'd8025:data <=32'h0080FFBB;14'd8026:data <=32'h006DFFAA;14'd8027:data <=32'h0056FFA2;
14'd8028:data <=32'h003FFFA0;14'd8029:data <=32'h002EFFA5;14'd8030:data <=32'h0023FFAD;
14'd8031:data <=32'h001BFFB4;14'd8032:data <=32'h0018FFBB;14'd8033:data <=32'h0015FFBD;
14'd8034:data <=32'h0011FFBC;14'd8035:data <=32'h000BFFBE;14'd8036:data <=32'h0003FFC2;
14'd8037:data <=32'hFFFBFFC8;14'd8038:data <=32'hFFF7FFD2;14'd8039:data <=32'hFFF8FFDF;
14'd8040:data <=32'hFFFEFFEA;14'd8041:data <=32'h0009FFF3;14'd8042:data <=32'h0018FFF5;
14'd8043:data <=32'h0028FFF3;14'd8044:data <=32'h0038FFEA;14'd8045:data <=32'h0045FFDD;
14'd8046:data <=32'h0051FFCA;14'd8047:data <=32'h0058FFB4;14'd8048:data <=32'h005BFF98;
14'd8049:data <=32'h0058FF77;14'd8050:data <=32'h004BFF54;14'd8051:data <=32'h0033FF2F;
14'd8052:data <=32'h000DFF0E;14'd8053:data <=32'hFFDAFEF6;14'd8054:data <=32'hFF9BFEED;
14'd8055:data <=32'hFF58FEF6;14'd8056:data <=32'hFF19FF13;14'd8057:data <=32'hFEE2FF43;
14'd8058:data <=32'hFEBAFF80;14'd8059:data <=32'hFEA4FFC4;14'd8060:data <=32'hFEA0000A;
14'd8061:data <=32'hFEAB004D;14'd8062:data <=32'hFEC40088;14'd8063:data <=32'hFEE900BB;
14'd8064:data <=32'hFF3E0034;14'd8065:data <=32'hFF2D005C;14'd8066:data <=32'hFF170088;
14'd8067:data <=32'hFEFE00CE;14'd8068:data <=32'hFF6F00D9;14'd8069:data <=32'hFF9800DE;
14'd8070:data <=32'hFFBE00DA;14'd8071:data <=32'hFFDD00CF;14'd8072:data <=32'hFFF200C1;
14'd8073:data <=32'h000100B5;14'd8074:data <=32'h000B00AE;14'd8075:data <=32'h001700AB;
14'd8076:data <=32'h002700A8;14'd8077:data <=32'h003B00A5;14'd8078:data <=32'h0050009C;
14'd8079:data <=32'h0066008C;14'd8080:data <=32'h00760076;14'd8081:data <=32'h0080005E;
14'd8082:data <=32'h00830045;14'd8083:data <=32'h007F002F;14'd8084:data <=32'h0078001D;
14'd8085:data <=32'h0070000D;14'd8086:data <=32'h00670002;14'd8087:data <=32'h005DFFF7;
14'd8088:data <=32'h0050FFF0;14'd8089:data <=32'h0042FFEC;14'd8090:data <=32'h0035FFEC;
14'd8091:data <=32'h0028FFF3;14'd8092:data <=32'h0020FFFE;14'd8093:data <=32'h001F000B;
14'd8094:data <=32'h00270018;14'd8095:data <=32'h00350020;14'd8096:data <=32'h00460022;
14'd8097:data <=32'h00560017;14'd8098:data <=32'h00630007;14'd8099:data <=32'h0067FFF3;
14'd8100:data <=32'h0065FFDF;14'd8101:data <=32'h0059FFCF;14'd8102:data <=32'h004BFFC6;
14'd8103:data <=32'h003BFFC2;14'd8104:data <=32'h002DFFC5;14'd8105:data <=32'h0023FFCC;
14'd8106:data <=32'h0020FFD5;14'd8107:data <=32'h0020FFDD;14'd8108:data <=32'h0025FFE5;
14'd8109:data <=32'h002DFFEB;14'd8110:data <=32'h0038FFED;14'd8111:data <=32'h0046FFEB;
14'd8112:data <=32'h0057FFE3;14'd8113:data <=32'h0068FFD4;14'd8114:data <=32'h0076FFBB;
14'd8115:data <=32'h007EFF9C;14'd8116:data <=32'h007CFF76;14'd8117:data <=32'h006CFF4D;
14'd8118:data <=32'h004EFF27;14'd8119:data <=32'h0023FF0D;14'd8120:data <=32'hFFF2FEFF;
14'd8121:data <=32'hFFBEFEFF;14'd8122:data <=32'hFF8DFF0D;14'd8123:data <=32'hFF63FF25;
14'd8124:data <=32'hFF43FF43;14'd8125:data <=32'hFF29FF65;14'd8126:data <=32'hFF18FF88;
14'd8127:data <=32'hFF0CFFAA;14'd8128:data <=32'hFEE4FF8E;14'd8129:data <=32'hFEBCFFBF;
14'd8130:data <=32'hFEAFFFE8;14'd8131:data <=32'hFEF5FFB4;14'd8132:data <=32'hFF2FFFC9;
14'd8133:data <=32'hFF26FFE1;14'd8134:data <=32'hFF1FFFF9;14'd8135:data <=32'hFF1A0015;
14'd8136:data <=32'hFF150032;14'd8137:data <=32'hFF130054;14'd8138:data <=32'hFF18007C;
14'd8139:data <=32'hFF2600A8;14'd8140:data <=32'hFF4200D3;14'd8141:data <=32'hFF6D00F7;
14'd8142:data <=32'hFFA00111;14'd8143:data <=32'hFFDC011A;14'd8144:data <=32'h00160111;
14'd8145:data <=32'h004900FB;14'd8146:data <=32'h007300D8;14'd8147:data <=32'h008F00B0;
14'd8148:data <=32'h00A00085;14'd8149:data <=32'h00A50059;14'd8150:data <=32'h00A00032;
14'd8151:data <=32'h0093000E;14'd8152:data <=32'h007FFFF0;14'd8153:data <=32'h0063FFD9;
14'd8154:data <=32'h0044FFCE;14'd8155:data <=32'h0023FFCC;14'd8156:data <=32'h0004FFD6;
14'd8157:data <=32'hFFECFFEB;14'd8158:data <=32'hFFE00007;14'd8159:data <=32'hFFE00023;
14'd8160:data <=32'hFFEA003D;14'd8161:data <=32'hFFFD004E;14'd8162:data <=32'h00140057;
14'd8163:data <=32'h00290057;14'd8164:data <=32'h003C0051;14'd8165:data <=32'h00490047;
14'd8166:data <=32'h0051003D;14'd8167:data <=32'h00590035;14'd8168:data <=32'h005F002D;
14'd8169:data <=32'h00650027;14'd8170:data <=32'h006C001F;14'd8171:data <=32'h00740015;
14'd8172:data <=32'h007B000A;14'd8173:data <=32'h007FFFFC;14'd8174:data <=32'h0082FFEE;
14'd8175:data <=32'h0082FFE0;14'd8176:data <=32'h0083FFD2;14'd8177:data <=32'h0082FFC5;
14'd8178:data <=32'h0082FFB5;14'd8179:data <=32'h007FFFA2;14'd8180:data <=32'h0078FF8D;
14'd8181:data <=32'h006CFF77;14'd8182:data <=32'h0058FF64;14'd8183:data <=32'h003FFF54;
14'd8184:data <=32'h0023FF4E;14'd8185:data <=32'h0005FF52;14'd8186:data <=32'hFFEFFF5B;
14'd8187:data <=32'hFFDEFF6A;14'd8188:data <=32'hFFD6FF78;14'd8189:data <=32'hFFD4FF82;
14'd8190:data <=32'hFFD5FF85;14'd8191:data <=32'hFFD4FF83;14'd8192:data <=32'hFF98FEE0;
14'd8193:data <=32'hFF56FEE6;14'd8194:data <=32'hFF2EFF0F;14'd8195:data <=32'hFFAFFF6B;
14'd8196:data <=32'hFFE2FF5B;14'd8197:data <=32'hFFC9FF4C;14'd8198:data <=32'hFFA8FF44;
14'd8199:data <=32'hFF82FF44;14'd8200:data <=32'hFF58FF4C;14'd8201:data <=32'hFF2AFF60;
14'd8202:data <=32'hFF00FF83;14'd8203:data <=32'hFEDFFFB5;14'd8204:data <=32'hFECBFFF2;
14'd8205:data <=32'hFECB0034;14'd8206:data <=32'hFEDD0074;14'd8207:data <=32'hFF0300AC;
14'd8208:data <=32'hFF3200D6;14'd8209:data <=32'hFF6900EF;14'd8210:data <=32'hFFA100F8;
14'd8211:data <=32'hFFD400F5;14'd8212:data <=32'h000200E7;14'd8213:data <=32'h002900D2;
14'd8214:data <=32'h004800B7;14'd8215:data <=32'h00600096;14'd8216:data <=32'h006F0073;
14'd8217:data <=32'h0075004E;14'd8218:data <=32'h0070002A;14'd8219:data <=32'h005F000C;
14'd8220:data <=32'h004AFFF7;14'd8221:data <=32'h002FFFEB;14'd8222:data <=32'h0016FFEA;
14'd8223:data <=32'h0001FFEF;14'd8224:data <=32'hFFF3FFFA;14'd8225:data <=32'hFFE60007;
14'd8226:data <=32'hFFE10013;14'd8227:data <=32'hFFDE001F;14'd8228:data <=32'hFFDA002A;
14'd8229:data <=32'hFFD70036;14'd8230:data <=32'hFFD70047;14'd8231:data <=32'hFFD8005C;
14'd8232:data <=32'hFFE10072;14'd8233:data <=32'hFFF30089;14'd8234:data <=32'h000D009B;
14'd8235:data <=32'h002E00A7;14'd8236:data <=32'h005300A9;14'd8237:data <=32'h007A00A0;
14'd8238:data <=32'h009D008F;14'd8239:data <=32'h00BC0075;14'd8240:data <=32'h00D30054;
14'd8241:data <=32'h00E5002F;14'd8242:data <=32'h00EE0007;14'd8243:data <=32'h00EFFFDC;
14'd8244:data <=32'h00E7FFB1;14'd8245:data <=32'h00D5FF88;14'd8246:data <=32'h00B8FF64;
14'd8247:data <=32'h0092FF48;14'd8248:data <=32'h0064FF3A;14'd8249:data <=32'h0039FF3A;
14'd8250:data <=32'h0011FF48;14'd8251:data <=32'hFFF5FF61;14'd8252:data <=32'hFFE7FF7D;
14'd8253:data <=32'hFFE5FF98;14'd8254:data <=32'hFFEFFFAB;14'd8255:data <=32'hFFFEFFB5;
14'd8256:data <=32'h0057FF4F;14'd8257:data <=32'h0040FF2D;14'd8258:data <=32'h0011FF24;
14'd8259:data <=32'hFFDFFF86;14'd8260:data <=32'h0021FF7D;14'd8261:data <=32'h0019FF6D;
14'd8262:data <=32'h000BFF5E;14'd8263:data <=32'hFFF7FF4F;14'd8264:data <=32'hFFDDFF43;
14'd8265:data <=32'hFFBBFF3D;14'd8266:data <=32'hFF95FF40;14'd8267:data <=32'hFF6DFF4F;
14'd8268:data <=32'hFF4AFF6B;14'd8269:data <=32'hFF30FF8F;14'd8270:data <=32'hFF22FFBB;
14'd8271:data <=32'hFF22FFE6;14'd8272:data <=32'hFF2C000B;14'd8273:data <=32'hFF3E002A;
14'd8274:data <=32'hFF520041;14'd8275:data <=32'hFF650050;14'd8276:data <=32'hFF78005C;
14'd8277:data <=32'hFF890067;14'd8278:data <=32'hFF9B0070;14'd8279:data <=32'hFFAE0077;
14'd8280:data <=32'hFFC3007B;14'd8281:data <=32'hFFD7007A;14'd8282:data <=32'hFFEC0074;
14'd8283:data <=32'hFFFC006A;14'd8284:data <=32'h0007005D;14'd8285:data <=32'h00110052;
14'd8286:data <=32'h00150046;14'd8287:data <=32'h0019003C;14'd8288:data <=32'h001D002F;
14'd8289:data <=32'h001E0023;14'd8290:data <=32'h001D0013;14'd8291:data <=32'h00160003;
14'd8292:data <=32'h0007FFF3;14'd8293:data <=32'hFFF0FFE9;14'd8294:data <=32'hFFD4FFE8;
14'd8295:data <=32'hFFB7FFF3;14'd8296:data <=32'hFF9D000A;14'd8297:data <=32'hFF8B002C;
14'd8298:data <=32'hFF850054;14'd8299:data <=32'hFF8C007E;14'd8300:data <=32'hFFA200A6;
14'd8301:data <=32'hFFC300C6;14'd8302:data <=32'hFFEC00DC;14'd8303:data <=32'h001800E8;
14'd8304:data <=32'h004700E9;14'd8305:data <=32'h007600E0;14'd8306:data <=32'h00A200CC;
14'd8307:data <=32'h00C900AE;14'd8308:data <=32'h00EB0088;14'd8309:data <=32'h01010059;
14'd8310:data <=32'h010A0027;14'd8311:data <=32'h0106FFF2;14'd8312:data <=32'h00F4FFC5;
14'd8313:data <=32'h00D8FFA1;14'd8314:data <=32'h00B7FF8A;14'd8315:data <=32'h0095FF80;
14'd8316:data <=32'h007CFF7E;14'd8317:data <=32'h0069FF82;14'd8318:data <=32'h005EFF86;
14'd8319:data <=32'h0058FF87;14'd8320:data <=32'h0039FFBC;14'd8321:data <=32'h0047FFB5;
14'd8322:data <=32'h004BFF9A;14'd8323:data <=32'h0040FF3F;14'd8324:data <=32'h0068FF35;
14'd8325:data <=32'h0049FF29;14'd8326:data <=32'h0029FF23;14'd8327:data <=32'h0007FF24;
14'd8328:data <=32'hFFE9FF29;14'd8329:data <=32'hFFC9FF31;14'd8330:data <=32'hFFADFF40;
14'd8331:data <=32'hFF90FF56;14'd8332:data <=32'hFF7AFF73;14'd8333:data <=32'hFF6EFF95;
14'd8334:data <=32'hFF6CFFB8;14'd8335:data <=32'hFF75FFD7;14'd8336:data <=32'hFF87FFEE;
14'd8337:data <=32'hFF9DFFF9;14'd8338:data <=32'hFFB1FFFB;14'd8339:data <=32'hFFBEFFF4;
14'd8340:data <=32'hFFC3FFE9;14'd8341:data <=32'hFFC0FFE1;14'd8342:data <=32'hFFB7FFDC;
14'd8343:data <=32'hFFACFFDD;14'd8344:data <=32'hFFA2FFE4;14'd8345:data <=32'hFF99FFEF;
14'd8346:data <=32'hFF95FFFB;14'd8347:data <=32'hFF92000A;14'd8348:data <=32'hFF930019;
14'd8349:data <=32'hFF970028;14'd8350:data <=32'hFF9E0038;14'd8351:data <=32'hFFAA0047;
14'd8352:data <=32'hFFBC0051;14'd8353:data <=32'hFFD20056;14'd8354:data <=32'hFFE90051;
14'd8355:data <=32'hFFFC0045;14'd8356:data <=32'h00090032;14'd8357:data <=32'h000C001A;
14'd8358:data <=32'h00040003;14'd8359:data <=32'hFFF2FFF2;14'd8360:data <=32'hFFDAFFE9;
14'd8361:data <=32'hFFBFFFEC;14'd8362:data <=32'hFFA7FFFA;14'd8363:data <=32'hFF96000F;
14'd8364:data <=32'hFF8B0029;14'd8365:data <=32'hFF890046;14'd8366:data <=32'hFF8E0061;
14'd8367:data <=32'hFF97007A;14'd8368:data <=32'hFFA60092;14'd8369:data <=32'hFFB900A7;
14'd8370:data <=32'hFFD000B8;14'd8371:data <=32'hFFEC00C7;14'd8372:data <=32'h000C00CF;
14'd8373:data <=32'h002D00D0;14'd8374:data <=32'h004E00C9;14'd8375:data <=32'h006B00BD;
14'd8376:data <=32'h008400AD;14'd8377:data <=32'h0098009A;14'd8378:data <=32'h00A80089;
14'd8379:data <=32'h00B7007A;14'd8380:data <=32'h00C9006A;14'd8381:data <=32'h00DC0057;
14'd8382:data <=32'h00F3003E;14'd8383:data <=32'h0107001D;14'd8384:data <=32'h005BFFB9;
14'd8385:data <=32'h005EFFC0;14'd8386:data <=32'h0074FFC8;14'd8387:data <=32'h0112FFBB;
14'd8388:data <=32'h0144FF84;14'd8389:data <=32'h0123FF49;14'd8390:data <=32'h00F6FF1A;
14'd8391:data <=32'h00C1FEF7;14'd8392:data <=32'h0088FEE1;14'd8393:data <=32'h004DFED8;
14'd8394:data <=32'h0011FEDB;14'd8395:data <=32'hFFD9FEED;14'd8396:data <=32'hFFA6FF0B;
14'd8397:data <=32'hFF80FF37;14'd8398:data <=32'hFF6AFF69;14'd8399:data <=32'hFF66FF9D;
14'd8400:data <=32'hFF71FFCB;14'd8401:data <=32'hFF89FFED;14'd8402:data <=32'hFFA80000;
14'd8403:data <=32'hFFC50006;14'd8404:data <=32'hFFDE0000;14'd8405:data <=32'hFFEEFFF3;
14'd8406:data <=32'hFFF5FFE4;14'd8407:data <=32'hFFF5FFD7;14'd8408:data <=32'hFFF1FFCC;
14'd8409:data <=32'hFFE9FFC4;14'd8410:data <=32'hFFE1FFBE;14'd8411:data <=32'hFFD7FFBB;
14'd8412:data <=32'hFFC9FFBA;14'd8413:data <=32'hFFBCFFBD;14'd8414:data <=32'hFFAFFFC4;
14'd8415:data <=32'hFFA4FFD0;14'd8416:data <=32'hFF9EFFE0;14'd8417:data <=32'hFF9DFFF0;
14'd8418:data <=32'hFFA1FFFF;14'd8419:data <=32'hFFAA0009;14'd8420:data <=32'hFFB4000D;
14'd8421:data <=32'hFFBB000C;14'd8422:data <=32'hFFBE0009;14'd8423:data <=32'hFFBC0006;
14'd8424:data <=32'hFFB60005;14'd8425:data <=32'hFFAF0009;14'd8426:data <=32'hFFAA0012;
14'd8427:data <=32'hFFA8001D;14'd8428:data <=32'hFFAC0027;14'd8429:data <=32'hFFB20031;
14'd8430:data <=32'hFFB90035;14'd8431:data <=32'hFFBF0036;14'd8432:data <=32'hFFC10034;
14'd8433:data <=32'hFFBF0032;14'd8434:data <=32'hFFB90033;14'd8435:data <=32'hFFB20038;
14'd8436:data <=32'hFFAA0042;14'd8437:data <=32'hFFA40050;14'd8438:data <=32'hFFA20062;
14'd8439:data <=32'hFFA10076;14'd8440:data <=32'hFFA4008C;14'd8441:data <=32'hFFAC00A6;
14'd8442:data <=32'hFFB900C3;14'd8443:data <=32'hFFD000E3;14'd8444:data <=32'hFFF20100;
14'd8445:data <=32'h00210118;14'd8446:data <=32'h005B0125;14'd8447:data <=32'h009E0122;
14'd8448:data <=32'h008B0059;14'd8449:data <=32'h00A10059;14'd8450:data <=32'h00A90066;
14'd8451:data <=32'h00D700D0;14'd8452:data <=32'h014100A0;14'd8453:data <=32'h0156005D;
14'd8454:data <=32'h015C001B;14'd8455:data <=32'h0150FFDA;14'd8456:data <=32'h013BFFA0;
14'd8457:data <=32'h011BFF6C;14'd8458:data <=32'h00F1FF41;14'd8459:data <=32'h00BEFF22;
14'd8460:data <=32'h0087FF11;14'd8461:data <=32'h0051FF11;14'd8462:data <=32'h001FFF1D;
14'd8463:data <=32'hFFF8FF35;14'd8464:data <=32'hFFDDFF53;14'd8465:data <=32'hFFCFFF71;
14'd8466:data <=32'hFFCBFF8B;14'd8467:data <=32'hFFCCFF9E;14'd8468:data <=32'hFFCFFFAC;
14'd8469:data <=32'hFFD0FFB5;14'd8470:data <=32'hFFD1FFBD;14'd8471:data <=32'hFFD0FFC6;
14'd8472:data <=32'hFFD1FFD0;14'd8473:data <=32'hFFD6FFDB;14'd8474:data <=32'hFFDDFFE2;
14'd8475:data <=32'hFFE7FFE7;14'd8476:data <=32'hFFF0FFE7;14'd8477:data <=32'hFFFAFFE3;
14'd8478:data <=32'h0000FFDC;14'd8479:data <=32'h0001FFD3;14'd8480:data <=32'h0001FFCB;
14'd8481:data <=32'hFFFFFFC3;14'd8482:data <=32'hFFFAFFBB;14'd8483:data <=32'hFFF5FFB2;
14'd8484:data <=32'hFFECFFA9;14'd8485:data <=32'hFFDFFFA0;14'd8486:data <=32'hFFCEFF99;
14'd8487:data <=32'hFFB6FF97;14'd8488:data <=32'hFF9DFF9D;14'd8489:data <=32'hFF86FFAB;
14'd8490:data <=32'hFF72FFC2;14'd8491:data <=32'hFF68FFDE;14'd8492:data <=32'hFF67FFFD;
14'd8493:data <=32'hFF710019;14'd8494:data <=32'hFF82002F;14'd8495:data <=32'hFF980039;
14'd8496:data <=32'hFFAC003C;14'd8497:data <=32'hFFBD0036;14'd8498:data <=32'hFFC6002D;
14'd8499:data <=32'hFFC80022;14'd8500:data <=32'hFFC50018;14'd8501:data <=32'hFFBC0011;
14'd8502:data <=32'hFFAF000F;14'd8503:data <=32'hFF9F0011;14'd8504:data <=32'hFF8C0019;
14'd8505:data <=32'hFF79002A;14'd8506:data <=32'hFF690042;14'd8507:data <=32'hFF5C0066;
14'd8508:data <=32'hFF5B0091;14'd8509:data <=32'hFF6800C1;14'd8510:data <=32'hFF8500F0;
14'd8511:data <=32'hFFB30117;14'd8512:data <=32'hFFBC00D6;14'd8513:data <=32'hFFE10103;
14'd8514:data <=32'hFFFE0111;14'd8515:data <=32'hFFFC00ED;14'd8516:data <=32'h006600EA;
14'd8517:data <=32'h008600D1;14'd8518:data <=32'h009E00B8;14'd8519:data <=32'h00B0009B;
14'd8520:data <=32'h00BF0081;14'd8521:data <=32'h00CB0064;14'd8522:data <=32'h00D20045;
14'd8523:data <=32'h00D40026;14'd8524:data <=32'h00D00008;14'd8525:data <=32'h00C7FFED;
14'd8526:data <=32'h00B9FFD8;14'd8527:data <=32'h00AEFFC8;14'd8528:data <=32'h00A3FFBA;
14'd8529:data <=32'h0099FFAB;14'd8530:data <=32'h0090FF9D;14'd8531:data <=32'h0085FF8A;
14'd8532:data <=32'h0075FF76;14'd8533:data <=32'h005CFF65;14'd8534:data <=32'h003DFF59;
14'd8535:data <=32'h0018FF57;14'd8536:data <=32'hFFF5FF60;14'd8537:data <=32'hFFD8FF74;
14'd8538:data <=32'hFFC4FF90;14'd8539:data <=32'hFFBAFFAE;14'd8540:data <=32'hFFB9FFCB;
14'd8541:data <=32'hFFC1FFE5;14'd8542:data <=32'hFFD0FFF8;14'd8543:data <=32'hFFE30005;
14'd8544:data <=32'hFFF7000D;14'd8545:data <=32'h000F000D;14'd8546:data <=32'h00240007;
14'd8547:data <=32'h0039FFFA;14'd8548:data <=32'h0047FFE4;14'd8549:data <=32'h004FFFC8;
14'd8550:data <=32'h004EFFA9;14'd8551:data <=32'h0040FF89;14'd8552:data <=32'h0029FF71;
14'd8553:data <=32'h0009FF5F;14'd8554:data <=32'hFFE5FF5A;14'd8555:data <=32'hFFC3FF5F;
14'd8556:data <=32'hFFA6FF6F;14'd8557:data <=32'hFF91FF85;14'd8558:data <=32'hFF85FF9C;
14'd8559:data <=32'hFF80FFB0;14'd8560:data <=32'hFF7EFFC1;14'd8561:data <=32'hFF7FFFCC;
14'd8562:data <=32'hFF7EFFD6;14'd8563:data <=32'hFF7CFFDF;14'd8564:data <=32'hFF78FFE7;
14'd8565:data <=32'hFF72FFF2;14'd8566:data <=32'hFF6FFFFD;14'd8567:data <=32'hFF6C0009;
14'd8568:data <=32'hFF680016;14'd8569:data <=32'hFF650024;14'd8570:data <=32'hFF600033;
14'd8571:data <=32'hFF5C0047;14'd8572:data <=32'hFF5B0060;14'd8573:data <=32'hFF60007E;
14'd8574:data <=32'hFF70009D;14'd8575:data <=32'hFF8800B8;14'd8576:data <=32'hFF120034;
14'd8577:data <=32'hFF04007F;14'd8578:data <=32'hFF2100BC;14'd8579:data <=32'hFFCB00A6;
14'd8580:data <=32'h002200A2;14'd8581:data <=32'h002C008B;14'd8582:data <=32'h002E0077;
14'd8583:data <=32'h00280069;14'd8584:data <=32'h00230064;14'd8585:data <=32'h001E0065;
14'd8586:data <=32'h001F006A;14'd8587:data <=32'h00230071;14'd8588:data <=32'h002A0077;
14'd8589:data <=32'h0037007E;14'd8590:data <=32'h00460082;14'd8591:data <=32'h005A0086;
14'd8592:data <=32'h00730084;14'd8593:data <=32'h0090007D;14'd8594:data <=32'h00AE006A;
14'd8595:data <=32'h00C9004D;14'd8596:data <=32'h00DC0025;14'd8597:data <=32'h00E2FFF6;
14'd8598:data <=32'h00D8FFC5;14'd8599:data <=32'h00C0FF9B;14'd8600:data <=32'h009DFF7B;
14'd8601:data <=32'h0074FF68;14'd8602:data <=32'h004BFF64;14'd8603:data <=32'h0025FF69;
14'd8604:data <=32'h0006FF79;14'd8605:data <=32'hFFEEFF8E;14'd8606:data <=32'hFFDEFFA6;
14'd8607:data <=32'hFFD6FFBE;14'd8608:data <=32'hFFD4FFD7;14'd8609:data <=32'hFFD9FFEF;
14'd8610:data <=32'hFFE50004;14'd8611:data <=32'hFFF90014;14'd8612:data <=32'h000F001D;
14'd8613:data <=32'h0029001C;14'd8614:data <=32'h00410013;14'd8615:data <=32'h00540002;
14'd8616:data <=32'h0061FFEA;14'd8617:data <=32'h0066FFD1;14'd8618:data <=32'h0063FFBA;
14'd8619:data <=32'h005CFFA5;14'd8620:data <=32'h0051FF94;14'd8621:data <=32'h0047FF86;
14'd8622:data <=32'h003CFF78;14'd8623:data <=32'h0031FF68;14'd8624:data <=32'h0022FF57;
14'd8625:data <=32'h000EFF44;14'd8626:data <=32'hFFF1FF33;14'd8627:data <=32'hFFCEFF28;
14'd8628:data <=32'hFFA5FF24;14'd8629:data <=32'hFF79FF2E;14'd8630:data <=32'hFF50FF41;
14'd8631:data <=32'hFF2BFF5E;14'd8632:data <=32'hFF0FFF82;14'd8633:data <=32'hFEF9FFAB;
14'd8634:data <=32'hFEEBFFD9;14'd8635:data <=32'hFEE60008;14'd8636:data <=32'hFEEA0038;
14'd8637:data <=32'hFEF9006A;14'd8638:data <=32'hFF130097;14'd8639:data <=32'hFF3900BF;
14'd8640:data <=32'hFF54FFB6;14'd8641:data <=32'hFF26FFDC;14'd8642:data <=32'hFF0C0022;
14'd8643:data <=32'hFF7500C5;14'd8644:data <=32'hFFE400C8;14'd8645:data <=32'h000200AC;
14'd8646:data <=32'h0013008D;14'd8647:data <=32'h00160070;14'd8648:data <=32'h0012005C;
14'd8649:data <=32'h0009004E;14'd8650:data <=32'hFFFF0049;14'd8651:data <=32'hFFF60049;
14'd8652:data <=32'hFFEE004E;14'd8653:data <=32'hFFE80058;14'd8654:data <=32'hFFE70065;
14'd8655:data <=32'hFFEB0075;14'd8656:data <=32'hFFF70087;14'd8657:data <=32'h000B0096;
14'd8658:data <=32'h002600A1;14'd8659:data <=32'h004800A1;14'd8660:data <=32'h006A0096;
14'd8661:data <=32'h0087007F;14'd8662:data <=32'h009B0060;14'd8663:data <=32'h00A5003E;
14'd8664:data <=32'h00A3001D;14'd8665:data <=32'h009A0001;14'd8666:data <=32'h008BFFEC;
14'd8667:data <=32'h007BFFDE;14'd8668:data <=32'h006BFFD3;14'd8669:data <=32'h005EFFCD;
14'd8670:data <=32'h0051FFC8;14'd8671:data <=32'h0043FFC4;14'd8672:data <=32'h0035FFC2;
14'd8673:data <=32'h0026FFC4;14'd8674:data <=32'h0019FFCB;14'd8675:data <=32'h000FFFD4;
14'd8676:data <=32'h0009FFE1;14'd8677:data <=32'h0008FFEE;14'd8678:data <=32'h000AFFFA;
14'd8679:data <=32'h00110004;14'd8680:data <=32'h0019000B;14'd8681:data <=32'h00230012;
14'd8682:data <=32'h002D0016;14'd8683:data <=32'h003C001A;14'd8684:data <=32'h004C001C;
14'd8685:data <=32'h00630019;14'd8686:data <=32'h007D000F;14'd8687:data <=32'h0098FFFC;
14'd8688:data <=32'h00AFFFDB;14'd8689:data <=32'h00C0FFAF;14'd8690:data <=32'h00C0FF7D;
14'd8691:data <=32'h00B3FF46;14'd8692:data <=32'h0093FF14;14'd8693:data <=32'h0066FEEB;
14'd8694:data <=32'h002EFECD;14'd8695:data <=32'hFFEFFEBF;14'd8696:data <=32'hFFAFFEC1;
14'd8697:data <=32'hFF72FED0;14'd8698:data <=32'hFF38FEEE;14'd8699:data <=32'hFF06FF16;
14'd8700:data <=32'hFEDBFF4A;14'd8701:data <=32'hFEC0FF87;14'd8702:data <=32'hFEB3FFC9;
14'd8703:data <=32'hFEB8000D;14'd8704:data <=32'hFF52FFB2;14'd8705:data <=32'hFF33FFC9;
14'd8706:data <=32'hFF0AFFE5;14'd8707:data <=32'hFED2002A;14'd8708:data <=32'hFF330059;
14'd8709:data <=32'hFF4E0066;14'd8710:data <=32'hFF66006C;14'd8711:data <=32'hFF76006F;
14'd8712:data <=32'hFF830074;14'd8713:data <=32'hFF8F007B;14'd8714:data <=32'hFF9C0084;
14'd8715:data <=32'hFFAC008A;14'd8716:data <=32'hFFBE008F;14'd8717:data <=32'hFFD00090;
14'd8718:data <=32'hFFDF0090;14'd8719:data <=32'hFFED008D;14'd8720:data <=32'hFFF9008B;
14'd8721:data <=32'h0007008B;14'd8722:data <=32'h00170087;14'd8723:data <=32'h00280081;
14'd8724:data <=32'h00390075;14'd8725:data <=32'h00460064;14'd8726:data <=32'h004D004F;
14'd8727:data <=32'h004C003C;14'd8728:data <=32'h0044002B;14'd8729:data <=32'h00370022;
14'd8730:data <=32'h002B0020;14'd8731:data <=32'h00210025;14'd8732:data <=32'h001F002E;
14'd8733:data <=32'h00230038;14'd8734:data <=32'h002D003D;14'd8735:data <=32'h0039003D;
14'd8736:data <=32'h00440038;14'd8737:data <=32'h004E002E;14'd8738:data <=32'h00520022;
14'd8739:data <=32'h00530015;14'd8740:data <=32'h0050000B;14'd8741:data <=32'h004C0002;
14'd8742:data <=32'h0046FFFA;14'd8743:data <=32'h003EFFF5;14'd8744:data <=32'h0035FFF2;
14'd8745:data <=32'h002AFFF3;14'd8746:data <=32'h0021FFFA;14'd8747:data <=32'h00190007;
14'd8748:data <=32'h00190017;14'd8749:data <=32'h0020002B;14'd8750:data <=32'h0033003D;
14'd8751:data <=32'h004E0048;14'd8752:data <=32'h00710048;14'd8753:data <=32'h0098003A;
14'd8754:data <=32'h00B9001E;14'd8755:data <=32'h00D1FFF7;14'd8756:data <=32'h00DDFFC7;
14'd8757:data <=32'h00DBFF95;14'd8758:data <=32'h00CBFF66;14'd8759:data <=32'h00B2FF3C;
14'd8760:data <=32'h008FFF1A;14'd8761:data <=32'h0066FEFE;14'd8762:data <=32'h003AFEED;
14'd8763:data <=32'h000BFEE3;14'd8764:data <=32'hFFDBFEE3;14'd8765:data <=32'hFFA9FEED;
14'd8766:data <=32'hFF7BFF02;14'd8767:data <=32'hFF55FF22;14'd8768:data <=32'hFF4BFF1E;
14'd8769:data <=32'hFF1CFF39;14'd8770:data <=32'hFF05FF50;14'd8771:data <=32'hFF49FF2B;
14'd8772:data <=32'hFF76FF51;14'd8773:data <=32'hFF5FFF5B;14'd8774:data <=32'hFF44FF67;
14'd8775:data <=32'hFF27FF7A;14'd8776:data <=32'hFF0BFF99;14'd8777:data <=32'hFEF4FFC2;
14'd8778:data <=32'hFEE8FFF3;14'd8779:data <=32'hFEE90028;14'd8780:data <=32'hFEF7005B;
14'd8781:data <=32'hFF120087;14'd8782:data <=32'hFF3500AA;14'd8783:data <=32'hFF5D00C4;
14'd8784:data <=32'hFF8700D4;14'd8785:data <=32'hFFB400DB;14'd8786:data <=32'hFFE000DA;
14'd8787:data <=32'h000B00CE;14'd8788:data <=32'h003100B8;14'd8789:data <=32'h004F0097;
14'd8790:data <=32'h00620070;14'd8791:data <=32'h00670047;14'd8792:data <=32'h005D0020;
14'd8793:data <=32'h00470003;14'd8794:data <=32'h002AFFF2;14'd8795:data <=32'h000CFFEF;
14'd8796:data <=32'hFFF1FFF7;14'd8797:data <=32'hFFE00007;14'd8798:data <=32'hFFD6001B;
14'd8799:data <=32'hFFD6002F;14'd8800:data <=32'hFFDB003F;14'd8801:data <=32'hFFE5004C;
14'd8802:data <=32'hFFF10056;14'd8803:data <=32'hFFFD005C;14'd8804:data <=32'h000A0060;
14'd8805:data <=32'h00170062;14'd8806:data <=32'h0024005F;14'd8807:data <=32'h0030005B;
14'd8808:data <=32'h003B0055;14'd8809:data <=32'h0042004C;14'd8810:data <=32'h00460042;
14'd8811:data <=32'h0047003C;14'd8812:data <=32'h0048003A;14'd8813:data <=32'h0048003B;
14'd8814:data <=32'h004E003E;14'd8815:data <=32'h00590042;14'd8816:data <=32'h00690042;
14'd8817:data <=32'h007D003C;14'd8818:data <=32'h0090002D;14'd8819:data <=32'h009F0018;
14'd8820:data <=32'h00A7FFFE;14'd8821:data <=32'h00A7FFE3;14'd8822:data <=32'h00A1FFCB;
14'd8823:data <=32'h0095FFB7;14'd8824:data <=32'h0089FFA9;14'd8825:data <=32'h007DFF9F;
14'd8826:data <=32'h0074FF96;14'd8827:data <=32'h006DFF8C;14'd8828:data <=32'h0065FF82;
14'd8829:data <=32'h005BFF76;14'd8830:data <=32'h004FFF6B;14'd8831:data <=32'h0043FF61;
14'd8832:data <=32'h002EFECE;14'd8833:data <=32'hFFF4FEBE;14'd8834:data <=32'hFFCCFED5;
14'd8835:data <=32'h0034FF48;14'd8836:data <=32'h006AFF44;14'd8837:data <=32'h0054FF1E;
14'd8838:data <=32'h0030FEFC;14'd8839:data <=32'h0000FEE1;14'd8840:data <=32'hFFC4FED6;
14'd8841:data <=32'hFF83FEDD;14'd8842:data <=32'hFF44FEF7;14'd8843:data <=32'hFF11FF22;
14'd8844:data <=32'hFEEBFF58;14'd8845:data <=32'hFED3FF94;14'd8846:data <=32'hFECDFFD1;
14'd8847:data <=32'hFED4000C;14'd8848:data <=32'hFEE60043;14'd8849:data <=32'hFF030073;
14'd8850:data <=32'hFF29009B;14'd8851:data <=32'hFF5700B8;14'd8852:data <=32'hFF8B00C8;
14'd8853:data <=32'hFFBF00C9;14'd8854:data <=32'hFFEF00BB;14'd8855:data <=32'h001600A1;
14'd8856:data <=32'h0030007F;14'd8857:data <=32'h003C005A;14'd8858:data <=32'h003B0039;
14'd8859:data <=32'h0031001D;14'd8860:data <=32'h0022000C;14'd8861:data <=32'h00120001;
14'd8862:data <=32'h0004FFFC;14'd8863:data <=32'hFFF6FFFA;14'd8864:data <=32'hFFEBFFFA;
14'd8865:data <=32'hFFDEFFFC;14'd8866:data <=32'hFFD1FFFE;14'd8867:data <=32'hFFC30006;
14'd8868:data <=32'hFFB50012;14'd8869:data <=32'hFFAC0023;14'd8870:data <=32'hFFA70038;
14'd8871:data <=32'hFFA8004F;14'd8872:data <=32'hFFAE0067;14'd8873:data <=32'hFFBA007C;
14'd8874:data <=32'hFFCB008F;14'd8875:data <=32'hFFDF009E;14'd8876:data <=32'hFFF600AB;
14'd8877:data <=32'h000F00B4;14'd8878:data <=32'h002E00B8;14'd8879:data <=32'h004F00BA;
14'd8880:data <=32'h007200B1;14'd8881:data <=32'h0095009F;14'd8882:data <=32'h00B50083;
14'd8883:data <=32'h00CB005E;14'd8884:data <=32'h00D60033;14'd8885:data <=32'h00D30008;
14'd8886:data <=32'h00C3FFE2;14'd8887:data <=32'h00ABFFC6;14'd8888:data <=32'h008FFFB6;
14'd8889:data <=32'h0074FFB0;14'd8890:data <=32'h005EFFB5;14'd8891:data <=32'h004FFFBD;
14'd8892:data <=32'h0048FFC9;14'd8893:data <=32'h0046FFD3;14'd8894:data <=32'h004CFFDA;
14'd8895:data <=32'h0054FFDD;14'd8896:data <=32'h00B9FF94;14'd8897:data <=32'h00B4FF71;
14'd8898:data <=32'h0092FF5E;14'd8899:data <=32'h0052FFB7;14'd8900:data <=32'h009FFFBE;
14'd8901:data <=32'h00A7FF9C;14'd8902:data <=32'h00A4FF74;14'd8903:data <=32'h0094FF49;
14'd8904:data <=32'h0075FF23;14'd8905:data <=32'h0048FF08;14'd8906:data <=32'h0016FEFB;
14'd8907:data <=32'hFFE4FEFC;14'd8908:data <=32'hFFB6FF0B;14'd8909:data <=32'hFF90FF20;
14'd8910:data <=32'hFF72FF3D;14'd8911:data <=32'hFF5AFF5B;14'd8912:data <=32'hFF48FF7C;
14'd8913:data <=32'hFF3DFF9E;14'd8914:data <=32'hFF37FFC1;14'd8915:data <=32'hFF39FFE5;
14'd8916:data <=32'hFF430006;14'd8917:data <=32'hFF540023;14'd8918:data <=32'hFF6A0038;
14'd8919:data <=32'hFF830045;14'd8920:data <=32'hFF9A004B;14'd8921:data <=32'hFFAC004B;
14'd8922:data <=32'hFFBB0049;14'd8923:data <=32'hFFC70048;14'd8924:data <=32'hFFD20047;
14'd8925:data <=32'hFFDE0047;14'd8926:data <=32'hFFEC0045;14'd8927:data <=32'hFFFB003D;
14'd8928:data <=32'h000A0030;14'd8929:data <=32'h0013001C;14'd8930:data <=32'h00140004;
14'd8931:data <=32'h000DFFED;14'd8932:data <=32'hFFFCFFD9;14'd8933:data <=32'hFFE2FFCB;
14'd8934:data <=32'hFFC4FFC9;14'd8935:data <=32'hFFA6FFCF;14'd8936:data <=32'hFF8BFFDF;
14'd8937:data <=32'hFF75FFF7;14'd8938:data <=32'hFF630015;14'd8939:data <=32'hFF5A0038;
14'd8940:data <=32'hFF59005F;14'd8941:data <=32'hFF600087;14'd8942:data <=32'hFF7300B0;
14'd8943:data <=32'hFF9100D5;14'd8944:data <=32'hFFBC00F2;14'd8945:data <=32'hFFED0104;
14'd8946:data <=32'h00240106;14'd8947:data <=32'h005900F9;14'd8948:data <=32'h008700DE;
14'd8949:data <=32'h00A900B8;14'd8950:data <=32'h00BD008D;14'd8951:data <=32'h00C30064;
14'd8952:data <=32'h00BE0040;14'd8953:data <=32'h00B40026;14'd8954:data <=32'h00A70012;
14'd8955:data <=32'h009B0005;14'd8956:data <=32'h0092FFFC;14'd8957:data <=32'h008AFFF6;
14'd8958:data <=32'h0084FFF0;14'd8959:data <=32'h0081FFED;14'd8960:data <=32'h0053000E;
14'd8961:data <=32'h00660015;14'd8962:data <=32'h00770005;14'd8963:data <=32'h0086FFB6;
14'd8964:data <=32'h00C1FFC2;14'd8965:data <=32'h00BDFFA6;14'd8966:data <=32'h00B2FF88;
14'd8967:data <=32'h009FFF6B;14'd8968:data <=32'h0083FF52;14'd8969:data <=32'h005FFF43;
14'd8970:data <=32'h003AFF3E;14'd8971:data <=32'h0017FF45;14'd8972:data <=32'hFFF8FF54;
14'd8973:data <=32'hFFE6FF68;14'd8974:data <=32'hFFDCFF7C;14'd8975:data <=32'hFFD8FF8C;
14'd8976:data <=32'hFFD9FF97;14'd8977:data <=32'hFFDAFF9E;14'd8978:data <=32'hFFD8FFA1;
14'd8979:data <=32'hFFD5FFA3;14'd8980:data <=32'hFFD0FFA6;14'd8981:data <=32'hFFCCFFA7;
14'd8982:data <=32'hFFC7FFA9;14'd8983:data <=32'hFFC1FFAA;14'd8984:data <=32'hFFB8FFAC;
14'd8985:data <=32'hFFACFFAE;14'd8986:data <=32'hFF9DFFB7;14'd8987:data <=32'hFF8EFFC5;
14'd8988:data <=32'hFF83FFD9;14'd8989:data <=32'hFF7EFFF3;14'd8990:data <=32'hFF84000E;
14'd8991:data <=32'hFF940027;14'd8992:data <=32'hFFAB0037;14'd8993:data <=32'hFFC7003E;
14'd8994:data <=32'hFFE10039;14'd8995:data <=32'hFFF80029;14'd8996:data <=32'h00050014;
14'd8997:data <=32'h0008FFFC;14'd8998:data <=32'h0002FFE5;14'd8999:data <=32'hFFF5FFD2;
14'd9000:data <=32'hFFE2FFC5;14'd9001:data <=32'hFFCBFFBD;14'd9002:data <=32'hFFB3FFBC;
14'd9003:data <=32'hFF98FFC2;14'd9004:data <=32'hFF7EFFCF;14'd9005:data <=32'hFF66FFE4;
14'd9006:data <=32'hFF530000;14'd9007:data <=32'hFF480023;14'd9008:data <=32'hFF460049;
14'd9009:data <=32'hFF4F0070;14'd9010:data <=32'hFF620093;14'd9011:data <=32'hFF7D00AE;
14'd9012:data <=32'hFF9C00C0;14'd9013:data <=32'hFFBA00CA;14'd9014:data <=32'hFFD500CD;
14'd9015:data <=32'hFFEF00CE;14'd9016:data <=32'h000200CE;14'd9017:data <=32'h001600D1;
14'd9018:data <=32'h002E00D4;14'd9019:data <=32'h004800D7;14'd9020:data <=32'h006900D4;
14'd9021:data <=32'h008A00CA;14'd9022:data <=32'h00AC00B8;14'd9023:data <=32'h00CA009F;
14'd9024:data <=32'h00420000;14'd9025:data <=32'h003B0016;14'd9026:data <=32'h004E0033;
14'd9027:data <=32'h00EF005D;14'd9028:data <=32'h013C004C;14'd9029:data <=32'h0142000F;
14'd9030:data <=32'h013AFFD1;14'd9031:data <=32'h0125FF98;14'd9032:data <=32'h00FFFF63;
14'd9033:data <=32'h00CDFF3C;14'd9034:data <=32'h0093FF27;14'd9035:data <=32'h0059FF24;
14'd9036:data <=32'h0025FF32;14'd9037:data <=32'hFFFEFF4D;14'd9038:data <=32'hFFE4FF6F;
14'd9039:data <=32'hFFDAFF90;14'd9040:data <=32'hFFD9FFAD;14'd9041:data <=32'hFFE1FFC3;
14'd9042:data <=32'hFFEDFFD2;14'd9043:data <=32'hFFFAFFDA;14'd9044:data <=32'h0008FFDD;
14'd9045:data <=32'h0013FFDA;14'd9046:data <=32'h001EFFD3;14'd9047:data <=32'h0025FFC6;
14'd9048:data <=32'h0027FFB6;14'd9049:data <=32'h0022FFA4;14'd9050:data <=32'h0014FF93;
14'd9051:data <=32'h0000FF88;14'd9052:data <=32'hFFE8FF86;14'd9053:data <=32'hFFCFFF8D;
14'd9054:data <=32'hFFBBFF9B;14'd9055:data <=32'hFFB0FFAF;14'd9056:data <=32'hFFACFFC4;
14'd9057:data <=32'hFFB0FFD5;14'd9058:data <=32'hFFB8FFE1;14'd9059:data <=32'hFFC2FFE7;
14'd9060:data <=32'hFFCAFFE8;14'd9061:data <=32'hFFCEFFE7;14'd9062:data <=32'hFFD0FFE3;
14'd9063:data <=32'hFFCFFFE1;14'd9064:data <=32'hFFCDFFE1;14'd9065:data <=32'hFFCCFFE1;
14'd9066:data <=32'hFFCAFFE0;14'd9067:data <=32'hFFC8FFDF;14'd9068:data <=32'hFFC6FFDB;
14'd9069:data <=32'hFFC0FFD9;14'd9070:data <=32'hFFB8FFD6;14'd9071:data <=32'hFFADFFD8;
14'd9072:data <=32'hFFA2FFDB;14'd9073:data <=32'hFF97FFE2;14'd9074:data <=32'hFF8DFFE9;
14'd9075:data <=32'hFF85FFF1;14'd9076:data <=32'hFF7BFFFA;14'd9077:data <=32'hFF6F0002;
14'd9078:data <=32'hFF61000F;14'd9079:data <=32'hFF4F0021;14'd9080:data <=32'hFF3D003C;
14'd9081:data <=32'hFF310063;14'd9082:data <=32'hFF2E0093;14'd9083:data <=32'hFF3A00C7;
14'd9084:data <=32'hFF5800FA;14'd9085:data <=32'hFF840126;14'd9086:data <=32'hFFBC0147;
14'd9087:data <=32'hFFFD0158;14'd9088:data <=32'h00340077;14'd9089:data <=32'h00370084;
14'd9090:data <=32'h002E00A2;14'd9091:data <=32'h003F0131;14'd9092:data <=32'h00B8013A;
14'd9093:data <=32'h00F0010E;14'd9094:data <=32'h011C00D5;14'd9095:data <=32'h01390094;
14'd9096:data <=32'h0143004F;14'd9097:data <=32'h013A000A;14'd9098:data <=32'h011FFFCE;
14'd9099:data <=32'h00F8FFA0;14'd9100:data <=32'h00CBFF84;14'd9101:data <=32'h009DFF76;
14'd9102:data <=32'h0077FF77;14'd9103:data <=32'h0058FF7D;14'd9104:data <=32'h0041FF87;
14'd9105:data <=32'h0031FF92;14'd9106:data <=32'h0023FF9C;14'd9107:data <=32'h0019FFA6;
14'd9108:data <=32'h0010FFB1;14'd9109:data <=32'h000BFFBC;14'd9110:data <=32'h000BFFC7;
14'd9111:data <=32'h000EFFCF;14'd9112:data <=32'h0013FFD3;14'd9113:data <=32'h0019FFD4;
14'd9114:data <=32'h001CFFD1;14'd9115:data <=32'h001DFFCD;14'd9116:data <=32'h001BFFC9;
14'd9117:data <=32'h0017FFC7;14'd9118:data <=32'h0013FFC8;14'd9119:data <=32'h0013FFCA;
14'd9120:data <=32'h0016FFCA;14'd9121:data <=32'h001BFFC7;14'd9122:data <=32'h0020FFC0;
14'd9123:data <=32'h0022FFB4;14'd9124:data <=32'h001CFFA4;14'd9125:data <=32'h0013FF94;
14'd9126:data <=32'h0000FF8A;14'd9127:data <=32'hFFEAFF86;14'd9128:data <=32'hFFD3FF88;
14'd9129:data <=32'hFFC0FF92;14'd9130:data <=32'hFFB0FFA2;14'd9131:data <=32'hFFA8FFB4;
14'd9132:data <=32'hFFA6FFC4;14'd9133:data <=32'hFFA9FFD3;14'd9134:data <=32'hFFAEFFDF;
14'd9135:data <=32'hFFB5FFE7;14'd9136:data <=32'hFFBDFFE9;14'd9137:data <=32'hFFC5FFE9;
14'd9138:data <=32'hFFCDFFE5;14'd9139:data <=32'hFFD3FFDB;14'd9140:data <=32'hFFD2FFCD;
14'd9141:data <=32'hFFCAFFBB;14'd9142:data <=32'hFFB8FFAA;14'd9143:data <=32'hFF9CFF9C;
14'd9144:data <=32'hFF75FF9B;14'd9145:data <=32'hFF4AFFA8;14'd9146:data <=32'hFF21FFC4;
14'd9147:data <=32'hFEFFFFF1;14'd9148:data <=32'hFEEC0028;14'd9149:data <=32'hFEE90066;
14'd9150:data <=32'hFEF900A2;14'd9151:data <=32'hFF1800DA;14'd9152:data <=32'hFF5B0090;
14'd9153:data <=32'hFF5D00BF;14'd9154:data <=32'hFF5F00DB;14'd9155:data <=32'hFF5100D2;
14'd9156:data <=32'hFFB3010D;14'd9157:data <=32'hFFE20113;14'd9158:data <=32'h00100110;
14'd9159:data <=32'h003C0103;14'd9160:data <=32'h006300EC;14'd9161:data <=32'h008000D0;
14'd9162:data <=32'h009300B0;14'd9163:data <=32'h009D0091;14'd9164:data <=32'h00A00078;
14'd9165:data <=32'h00A40064;14'd9166:data <=32'h00A70054;14'd9167:data <=32'h00AE0043;
14'd9168:data <=32'h00B6002F;14'd9169:data <=32'h00BB0017;14'd9170:data <=32'h00BCFFFA;
14'd9171:data <=32'h00B5FFDD;14'd9172:data <=32'h00A6FFC0;14'd9173:data <=32'h0090FFA9;
14'd9174:data <=32'h0076FF99;14'd9175:data <=32'h005AFF92;14'd9176:data <=32'h0040FF92;
14'd9177:data <=32'h0029FF95;14'd9178:data <=32'h0013FF9D;14'd9179:data <=32'h0002FFAA;
14'd9180:data <=32'hFFF3FFBA;14'd9181:data <=32'hFFE9FFCF;14'd9182:data <=32'hFFE7FFE6;
14'd9183:data <=32'hFFEEFFFE;14'd9184:data <=32'hFFFD0013;14'd9185:data <=32'h0015001F;
14'd9186:data <=32'h00310022;14'd9187:data <=32'h004F0018;14'd9188:data <=32'h00660003;
14'd9189:data <=32'h0074FFE7;14'd9190:data <=32'h0077FFC6;14'd9191:data <=32'h006EFFA8;
14'd9192:data <=32'h005EFF8E;14'd9193:data <=32'h0045FF7C;14'd9194:data <=32'h002EFF73;
14'd9195:data <=32'h0016FF6F;14'd9196:data <=32'h0002FF72;14'd9197:data <=32'hFFF0FF76;
14'd9198:data <=32'hFFE0FF7D;14'd9199:data <=32'hFFD3FF85;14'd9200:data <=32'hFFC9FF8F;
14'd9201:data <=32'hFFC2FF99;14'd9202:data <=32'hFFBEFFA1;14'd9203:data <=32'hFFBEFFA9;
14'd9204:data <=32'hFFBFFFAB;14'd9205:data <=32'hFFBFFFA9;14'd9206:data <=32'hFFBAFFA1;
14'd9207:data <=32'hFFAFFF98;14'd9208:data <=32'hFF9BFF91;14'd9209:data <=32'hFF80FF91;
14'd9210:data <=32'hFF62FF9C;14'd9211:data <=32'hFF45FFB1;14'd9212:data <=32'hFF2FFFD0;
14'd9213:data <=32'hFF23FFF5;14'd9214:data <=32'hFF21001B;14'd9215:data <=32'hFF2A003E;
14'd9216:data <=32'hFF04FFAC;14'd9217:data <=32'hFED0FFE2;14'd9218:data <=32'hFEC5001B;
14'd9219:data <=32'hFF52003E;14'd9220:data <=32'hFF96006D;14'd9221:data <=32'hFFA2006E;
14'd9222:data <=32'hFFAC006F;14'd9223:data <=32'hFFB40071;14'd9224:data <=32'hFFBA0072;
14'd9225:data <=32'hFFBE0073;14'd9226:data <=32'hFFBE0077;14'd9227:data <=32'hFFBF0080;
14'd9228:data <=32'hFFC10090;14'd9229:data <=32'hFFC900A6;14'd9230:data <=32'hFFDC00BE;
14'd9231:data <=32'hFFF800D2;14'd9232:data <=32'h002100DE;14'd9233:data <=32'h004E00DE;
14'd9234:data <=32'h007B00CE;14'd9235:data <=32'h00A400B1;14'd9236:data <=32'h00C1008A;
14'd9237:data <=32'h00D1005E;14'd9238:data <=32'h00D50030;14'd9239:data <=32'h00CE0006;
14'd9240:data <=32'h00BFFFE1;14'd9241:data <=32'h00A9FFC1;14'd9242:data <=32'h008BFFA9;
14'd9243:data <=32'h006AFF99;14'd9244:data <=32'h0047FF92;14'd9245:data <=32'h0023FF96;
14'd9246:data <=32'h0003FFA4;14'd9247:data <=32'hFFEAFFBC;14'd9248:data <=32'hFFDDFFDB;
14'd9249:data <=32'hFFDCFFFB;14'd9250:data <=32'hFFE60019;14'd9251:data <=32'hFFFB002F;
14'd9252:data <=32'h0014003A;14'd9253:data <=32'h0030003C;14'd9254:data <=32'h00470036;
14'd9255:data <=32'h005A002A;14'd9256:data <=32'h0068001B;14'd9257:data <=32'h0072000B;
14'd9258:data <=32'h0079FFFC;14'd9259:data <=32'h0081FFED;14'd9260:data <=32'h0087FFDA;
14'd9261:data <=32'h008BFFC6;14'd9262:data <=32'h008CFFAD;14'd9263:data <=32'h0088FF93;
14'd9264:data <=32'h007DFF79;14'd9265:data <=32'h006DFF5F;14'd9266:data <=32'h0058FF4A;
14'd9267:data <=32'h003EFF38;14'd9268:data <=32'h0022FF2A;14'd9269:data <=32'h0004FF21;
14'd9270:data <=32'hFFE4FF1A;14'd9271:data <=32'hFFC0FF19;14'd9272:data <=32'hFF99FF1D;
14'd9273:data <=32'hFF70FF2B;14'd9274:data <=32'hFF48FF45;14'd9275:data <=32'hFF26FF68;
14'd9276:data <=32'hFF0EFF96;14'd9277:data <=32'hFF05FFC9;14'd9278:data <=32'hFF0BFFFA;
14'd9279:data <=32'hFF1F0026;14'd9280:data <=32'hFF99FF40;14'd9281:data <=32'hFF57FF41;
14'd9282:data <=32'hFF1DFF6B;14'd9283:data <=32'hFF410028;14'd9284:data <=32'hFF920057;
14'd9285:data <=32'hFFA80051;14'd9286:data <=32'hFFB90046;14'd9287:data <=32'hFFC2003A;
14'd9288:data <=32'hFFC6002C;14'd9289:data <=32'hFFC2001F;14'd9290:data <=32'hFFB60015;
14'd9291:data <=32'hFFA50013;14'd9292:data <=32'hFF90001A;14'd9293:data <=32'hFF7D002E;
14'd9294:data <=32'hFF71004C;14'd9295:data <=32'hFF730071;14'd9296:data <=32'hFF820097;
14'd9297:data <=32'hFF9D00B6;14'd9298:data <=32'hFFC300CB;14'd9299:data <=32'hFFED00D2;
14'd9300:data <=32'h001500CF;14'd9301:data <=32'h003800C0;14'd9302:data <=32'h005500AD;
14'd9303:data <=32'h006C0095;14'd9304:data <=32'h007C007B;14'd9305:data <=32'h00870060;
14'd9306:data <=32'h008C0044;14'd9307:data <=32'h008B0028;14'd9308:data <=32'h0084000C;
14'd9309:data <=32'h0075FFF5;14'd9310:data <=32'h0061FFE3;14'd9311:data <=32'h004BFFDB;
14'd9312:data <=32'h0035FFDA;14'd9313:data <=32'h0022FFE0;14'd9314:data <=32'h0015FFE9;
14'd9315:data <=32'h000CFFF5;14'd9316:data <=32'h00090000;14'd9317:data <=32'h00080009;
14'd9318:data <=32'h00070011;14'd9319:data <=32'h0005001B;14'd9320:data <=32'h00050027;
14'd9321:data <=32'h00080035;14'd9322:data <=32'h00120048;14'd9323:data <=32'h0023005A;
14'd9324:data <=32'h003C0067;14'd9325:data <=32'h005E006E;14'd9326:data <=32'h00830069;
14'd9327:data <=32'h00A90058;14'd9328:data <=32'h00CD003B;14'd9329:data <=32'h00E70013;
14'd9330:data <=32'h00F9FFE5;14'd9331:data <=32'h00FEFFB2;14'd9332:data <=32'h00F9FF7E;
14'd9333:data <=32'h00E7FF4A;14'd9334:data <=32'h00CAFF18;14'd9335:data <=32'h00A1FEEC;
14'd9336:data <=32'h006CFEC9;14'd9337:data <=32'h002DFEB2;14'd9338:data <=32'hFFE8FEAC;
14'd9339:data <=32'hFFA1FEB9;14'd9340:data <=32'hFF63FEDA;14'd9341:data <=32'hFF30FF0A;
14'd9342:data <=32'hFF0FFF44;14'd9343:data <=32'hFF03FF7F;14'd9344:data <=32'hFFC4FF65;
14'd9345:data <=32'hFFA4FF59;14'd9346:data <=32'hFF71FF50;14'd9347:data <=32'hFF0FFF83;
14'd9348:data <=32'hFF48FFCE;14'd9349:data <=32'hFF50FFE1;14'd9350:data <=32'hFF5BFFF3;
14'd9351:data <=32'hFF630001;14'd9352:data <=32'hFF6E000B;14'd9353:data <=32'hFF780012;
14'd9354:data <=32'hFF7F0016;14'd9355:data <=32'hFF820018;14'd9356:data <=32'hFF80001D;
14'd9357:data <=32'hFF7C0026;14'd9358:data <=32'hFF7A0036;14'd9359:data <=32'hFF7B004A;
14'd9360:data <=32'hFF850060;14'd9361:data <=32'hFF970072;14'd9362:data <=32'hFFAE007E;
14'd9363:data <=32'hFFC70082;14'd9364:data <=32'hFFDE007E;14'd9365:data <=32'hFFEE0074;
14'd9366:data <=32'hFFF90069;14'd9367:data <=32'hFFFD005E;14'd9368:data <=32'h00000058;
14'd9369:data <=32'h00020055;14'd9370:data <=32'h00050055;14'd9371:data <=32'h00090055;
14'd9372:data <=32'h000F0053;14'd9373:data <=32'h00150050;14'd9374:data <=32'h001B004C;
14'd9375:data <=32'h001F0049;14'd9376:data <=32'h00230046;14'd9377:data <=32'h00280042;
14'd9378:data <=32'h002E003F;14'd9379:data <=32'h00350038;14'd9380:data <=32'h003A002E;
14'd9381:data <=32'h003B0020;14'd9382:data <=32'h00370013;14'd9383:data <=32'h002B0007;
14'd9384:data <=32'h00190001;14'd9385:data <=32'h00060004;14'd9386:data <=32'hFFF20011;
14'd9387:data <=32'hFFE60028;14'd9388:data <=32'hFFE30046;14'd9389:data <=32'hFFED0065;
14'd9390:data <=32'h00040081;14'd9391:data <=32'h00250095;14'd9392:data <=32'h004D009E;
14'd9393:data <=32'h0076009C;14'd9394:data <=32'h00A0008E;14'd9395:data <=32'h00C60076;
14'd9396:data <=32'h00E70055;14'd9397:data <=32'h0102002C;14'd9398:data <=32'h0112FFFC;
14'd9399:data <=32'h011AFFC7;14'd9400:data <=32'h0115FF8E;14'd9401:data <=32'h00FEFF57;
14'd9402:data <=32'h00DAFF27;14'd9403:data <=32'h00ABFF01;14'd9404:data <=32'h0076FEEC;
14'd9405:data <=32'h0040FEE5;14'd9406:data <=32'h000EFEEB;14'd9407:data <=32'hFFE6FEFB;
14'd9408:data <=32'hFFE4FF0F;14'd9409:data <=32'hFFC1FF0D;14'd9410:data <=32'hFFAEFF05;
14'd9411:data <=32'hFFE6FEE2;14'd9412:data <=32'hFFF6FF0D;14'd9413:data <=32'hFFD5FF09;
14'd9414:data <=32'hFFAEFF0E;14'd9415:data <=32'hFF86FF19;14'd9416:data <=32'hFF63FF2F;
14'd9417:data <=32'hFF45FF4A;14'd9418:data <=32'hFF2DFF6C;14'd9419:data <=32'hFF1AFF8E;
14'd9420:data <=32'hFF0EFFB6;14'd9421:data <=32'hFF07FFDF;14'd9422:data <=32'hFF09000B;
14'd9423:data <=32'hFF160039;14'd9424:data <=32'hFF2D0062;14'd9425:data <=32'hFF510084;
14'd9426:data <=32'hFF7D0099;14'd9427:data <=32'hFFAC009F;14'd9428:data <=32'hFFD70097;
14'd9429:data <=32'hFFF90082;14'd9430:data <=32'h00100064;14'd9431:data <=32'h00180047;
14'd9432:data <=32'h0017002B;14'd9433:data <=32'h000D0017;14'd9434:data <=32'hFFFF000A;
14'd9435:data <=32'hFFF00004;14'd9436:data <=32'hFFE10004;14'd9437:data <=32'hFFD30007;
14'd9438:data <=32'hFFC70011;14'd9439:data <=32'hFFBF001B;14'd9440:data <=32'hFFBA002A;
14'd9441:data <=32'hFFBA003A;14'd9442:data <=32'hFFC1004C;14'd9443:data <=32'hFFCE005A;
14'd9444:data <=32'hFFDE0062;14'd9445:data <=32'hFFF00065;14'd9446:data <=32'h00000060;
14'd9447:data <=32'h000C0055;14'd9448:data <=32'h0010004A;14'd9449:data <=32'h000D0041;
14'd9450:data <=32'h0006003D;14'd9451:data <=32'hFFFD0040;14'd9452:data <=32'hFFF7004A;
14'd9453:data <=32'hFFF70059;14'd9454:data <=32'hFFFE0067;14'd9455:data <=32'h000C0075;
14'd9456:data <=32'h0020007D;14'd9457:data <=32'h00340081;14'd9458:data <=32'h0048007F;
14'd9459:data <=32'h005B007A;14'd9460:data <=32'h006E0072;14'd9461:data <=32'h007E0068;
14'd9462:data <=32'h0091005B;14'd9463:data <=32'h00A0004A;14'd9464:data <=32'h00AE0036;
14'd9465:data <=32'h00B90020;14'd9466:data <=32'h00BC0006;14'd9467:data <=32'h00BBFFEE;
14'd9468:data <=32'h00B6FFD9;14'd9469:data <=32'h00AFFFC8;14'd9470:data <=32'h00ABFFBC;
14'd9471:data <=32'h00AAFFAE;14'd9472:data <=32'h00B2FF25;14'd9473:data <=32'h0093FF05;
14'd9474:data <=32'h007AFF05;14'd9475:data <=32'h00C3FF7D;14'd9476:data <=32'h00F1FF7E;
14'd9477:data <=32'h00E3FF48;14'd9478:data <=32'h00C5FF15;14'd9479:data <=32'h0098FEE9;
14'd9480:data <=32'h0062FECB;14'd9481:data <=32'h0027FEBC;14'd9482:data <=32'hFFEAFEB9;
14'd9483:data <=32'hFFACFEC3;14'd9484:data <=32'hFF73FED9;14'd9485:data <=32'hFF3EFEFE;
14'd9486:data <=32'hFF12FF2D;14'd9487:data <=32'hFEF4FF68;14'd9488:data <=32'hFEE6FFA8;
14'd9489:data <=32'hFEEBFFEA;14'd9490:data <=32'hFF020024;14'd9491:data <=32'hFF280052;
14'd9492:data <=32'hFF550070;14'd9493:data <=32'hFF85007D;14'd9494:data <=32'hFFB0007A;
14'd9495:data <=32'hFFD3006F;14'd9496:data <=32'hFFED005C;14'd9497:data <=32'hFFFD0048;
14'd9498:data <=32'h00070033;14'd9499:data <=32'h000C0020;14'd9500:data <=32'h000B000E;
14'd9501:data <=32'h0006FFFE;14'd9502:data <=32'hFFFEFFEF;14'd9503:data <=32'hFFF0FFE4;
14'd9504:data <=32'hFFDFFFDC;14'd9505:data <=32'hFFCEFFDC;14'd9506:data <=32'hFFBBFFE1;
14'd9507:data <=32'hFFACFFEB;14'd9508:data <=32'hFFA3FFF8;14'd9509:data <=32'hFF9C0007;
14'd9510:data <=32'hFF990015;14'd9511:data <=32'hFF960022;14'd9512:data <=32'hFF94002F;
14'd9513:data <=32'hFF92003E;14'd9514:data <=32'hFF91004F;14'd9515:data <=32'hFF910065;
14'd9516:data <=32'hFF9A007D;14'd9517:data <=32'hFFA90097;14'd9518:data <=32'hFFC000AC;
14'd9519:data <=32'hFFE100BB;14'd9520:data <=32'h000400C0;14'd9521:data <=32'h002700BB;
14'd9522:data <=32'h004500AC;14'd9523:data <=32'h005D0097;14'd9524:data <=32'h006C007E;
14'd9525:data <=32'h00740066;14'd9526:data <=32'h00740052;14'd9527:data <=32'h00720041;
14'd9528:data <=32'h006C0032;14'd9529:data <=32'h00650028;14'd9530:data <=32'h005C0022;
14'd9531:data <=32'h00530021;14'd9532:data <=32'h004C0027;14'd9533:data <=32'h004A0032;
14'd9534:data <=32'h004F0041;14'd9535:data <=32'h00610050;14'd9536:data <=32'h00D70018;
14'd9537:data <=32'h00ECFFFD;14'd9538:data <=32'h00E1FFE4;14'd9539:data <=32'h00940028;
14'd9540:data <=32'h00E20041;14'd9541:data <=32'h00FB0015;14'd9542:data <=32'h0107FFE3;
14'd9543:data <=32'h0105FFAD;14'd9544:data <=32'h00F4FF7C;14'd9545:data <=32'h00DBFF51;
14'd9546:data <=32'h00B9FF2C;14'd9547:data <=32'h0092FF0F;14'd9548:data <=32'h0065FEFA;
14'd9549:data <=32'h0032FEEF;14'd9550:data <=32'hFFFFFEEE;14'd9551:data <=32'hFFCBFEFB;
14'd9552:data <=32'hFFA0FF16;14'd9553:data <=32'hFF7EFF39;14'd9554:data <=32'hFF67FF62;
14'd9555:data <=32'hFF5FFF8B;14'd9556:data <=32'hFF61FFAE;14'd9557:data <=32'hFF6AFFCB;
14'd9558:data <=32'hFF75FFE0;14'd9559:data <=32'hFF81FFEF;14'd9560:data <=32'hFF8AFFFC;
14'd9561:data <=32'hFF940008;14'd9562:data <=32'hFF9D0015;14'd9563:data <=32'hFFAB0021;
14'd9564:data <=32'hFFBB002A;14'd9565:data <=32'hFFCE002E;14'd9566:data <=32'hFFE4002B;
14'd9567:data <=32'hFFF60022;14'd9568:data <=32'h00030013;14'd9569:data <=32'h000B0001;
14'd9570:data <=32'h000CFFED;14'd9571:data <=32'h0007FFDA;14'd9572:data <=32'hFFFDFFC8;
14'd9573:data <=32'hFFEFFFBA;14'd9574:data <=32'hFFDCFFAE;14'd9575:data <=32'hFFC5FFA6;
14'd9576:data <=32'hFFA8FFA2;14'd9577:data <=32'hFF88FFA8;14'd9578:data <=32'hFF66FFB7;
14'd9579:data <=32'hFF48FFD2;14'd9580:data <=32'hFF30FFF9;14'd9581:data <=32'hFF240027;
14'd9582:data <=32'hFF280059;14'd9583:data <=32'hFF390089;14'd9584:data <=32'hFF5800B2;
14'd9585:data <=32'hFF8100CE;14'd9586:data <=32'hFFAE00DD;14'd9587:data <=32'hFFD900E0;
14'd9588:data <=32'h000000D8;14'd9589:data <=32'h002000C9;14'd9590:data <=32'h003800B5;
14'd9591:data <=32'h004A00A0;14'd9592:data <=32'h0056008A;14'd9593:data <=32'h005D0076;
14'd9594:data <=32'h005E0063;14'd9595:data <=32'h00590053;14'd9596:data <=32'h00500049;
14'd9597:data <=32'h00460047;14'd9598:data <=32'h003F004D;14'd9599:data <=32'h003F005B;
14'd9600:data <=32'h001E0065;14'd9601:data <=32'h00350083;14'd9602:data <=32'h00550081;
14'd9603:data <=32'h007C003E;14'd9604:data <=32'h00BC005F;14'd9605:data <=32'h00CC003F;
14'd9606:data <=32'h00D4001D;14'd9607:data <=32'h00D2FFF8;14'd9608:data <=32'h00C7FFD8;
14'd9609:data <=32'h00B6FFC0;14'd9610:data <=32'h00A4FFAE;14'd9611:data <=32'h0092FF9F;
14'd9612:data <=32'h0081FF95;14'd9613:data <=32'h0070FF8C;14'd9614:data <=32'h005EFF85;
14'd9615:data <=32'h004DFF81;14'd9616:data <=32'h003BFF82;14'd9617:data <=32'h002DFF87;
14'd9618:data <=32'h0022FF8B;14'd9619:data <=32'h001DFF90;14'd9620:data <=32'h0019FF91;
14'd9621:data <=32'h0017FF8C;14'd9622:data <=32'h0010FF84;14'd9623:data <=32'h0003FF7B;
14'd9624:data <=32'hFFEFFF74;14'd9625:data <=32'hFFD6FF75;14'd9626:data <=32'hFFBCFF7F;
14'd9627:data <=32'hFFA5FF91;14'd9628:data <=32'hFF96FFAC;14'd9629:data <=32'hFF91FFC8;
14'd9630:data <=32'hFF96FFE4;14'd9631:data <=32'hFFA2FFFC;14'd9632:data <=32'hFFB5000B;
14'd9633:data <=32'hFFCA0015;14'd9634:data <=32'hFFE00016;14'd9635:data <=32'hFFF50013;
14'd9636:data <=32'h00060008;14'd9637:data <=32'h0015FFF8;14'd9638:data <=32'h001DFFE2;
14'd9639:data <=32'h0020FFC8;14'd9640:data <=32'h0018FFAB;14'd9641:data <=32'h0005FF91;
14'd9642:data <=32'hFFE9FF7D;14'd9643:data <=32'hFFC5FF72;14'd9644:data <=32'hFF9DFF72;
14'd9645:data <=32'hFF76FF81;14'd9646:data <=32'hFF55FF9C;14'd9647:data <=32'hFF3DFFBD;
14'd9648:data <=32'hFF31FFE4;14'd9649:data <=32'hFF2F0007;14'd9650:data <=32'hFF34002A;
14'd9651:data <=32'hFF3D0045;14'd9652:data <=32'hFF4A005C;14'd9653:data <=32'hFF560072;
14'd9654:data <=32'hFF640085;14'd9655:data <=32'hFF730099;14'd9656:data <=32'hFF8500AC;
14'd9657:data <=32'hFF9B00BC;14'd9658:data <=32'hFFB300C9;14'd9659:data <=32'hFFCD00D1;
14'd9660:data <=32'hFFE600D6;14'd9661:data <=32'hFFFF00D9;14'd9662:data <=32'h001700DB;
14'd9663:data <=32'h003100DB;14'd9664:data <=32'hFFEF001D;14'd9665:data <=32'hFFDB0043;
14'd9666:data <=32'hFFE80074;14'd9667:data <=32'h007E00CF;14'd9668:data <=32'h00D400E2;
14'd9669:data <=32'h00F500AE;14'd9670:data <=32'h01080073;14'd9671:data <=32'h01090037;
14'd9672:data <=32'h00F90002;14'd9673:data <=32'h00DDFFD8;14'd9674:data <=32'h00BBFFBA;
14'd9675:data <=32'h0098FFAA;14'd9676:data <=32'h0078FFA4;14'd9677:data <=32'h005BFFA5;
14'd9678:data <=32'h0043FFAD;14'd9679:data <=32'h0031FFB9;14'd9680:data <=32'h0024FFC8;
14'd9681:data <=32'h001FFFDA;14'd9682:data <=32'h0023FFEB;14'd9683:data <=32'h002EFFF8;
14'd9684:data <=32'h003FFFFE;14'd9685:data <=32'h0054FFFA;14'd9686:data <=32'h0065FFEA;
14'd9687:data <=32'h0070FFD3;14'd9688:data <=32'h006FFFB7;14'd9689:data <=32'h0064FF9C;
14'd9690:data <=32'h004FFF87;14'd9691:data <=32'h0034FF7B;14'd9692:data <=32'h0018FF79;
14'd9693:data <=32'h0000FF7F;14'd9694:data <=32'hFFEDFF8B;14'd9695:data <=32'hFFDFFF9A;
14'd9696:data <=32'hFFD8FFAA;14'd9697:data <=32'hFFD4FFB7;14'd9698:data <=32'hFFD3FFC4;
14'd9699:data <=32'hFFD6FFD0;14'd9700:data <=32'hFFDBFFDA;14'd9701:data <=32'hFFE3FFE3;
14'd9702:data <=32'hFFEDFFE7;14'd9703:data <=32'hFFFAFFE6;14'd9704:data <=32'h0003FFDF;
14'd9705:data <=32'h000CFFD4;14'd9706:data <=32'h000FFFC5;14'd9707:data <=32'h000AFFB5;
14'd9708:data <=32'h0000FFA7;14'd9709:data <=32'hFFF2FF9E;14'd9710:data <=32'hFFE4FF99;
14'd9711:data <=32'hFFD6FF98;14'd9712:data <=32'hFFCBFF98;14'd9713:data <=32'hFFC1FF97;
14'd9714:data <=32'hFFB6FF94;14'd9715:data <=32'hFFA6FF8F;14'd9716:data <=32'hFF91FF8A;
14'd9717:data <=32'hFF75FF8A;14'd9718:data <=32'hFF55FF91;14'd9719:data <=32'hFF32FFA5;
14'd9720:data <=32'hFF11FFC3;14'd9721:data <=32'hFEF8FFED;14'd9722:data <=32'hFEE9001C;
14'd9723:data <=32'hFEE40051;14'd9724:data <=32'hFEEC0085;14'd9725:data <=32'hFEFE00BA;
14'd9726:data <=32'hFF1B00EC;14'd9727:data <=32'hFF42011A;14'd9728:data <=32'hFFD30050;
14'd9729:data <=32'hFFBE0065;14'd9730:data <=32'hFFA5008F;14'd9731:data <=32'hFF900134;
14'd9732:data <=32'h00000171;14'd9733:data <=32'h004B015C;14'd9734:data <=32'h008B0136;
14'd9735:data <=32'h00BB0102;14'd9736:data <=32'h00D700C9;14'd9737:data <=32'h00E3008F;
14'd9738:data <=32'h00E0005D;14'd9739:data <=32'h00D30033;14'd9740:data <=32'h00C20010;
14'd9741:data <=32'h00ACFFF7;14'd9742:data <=32'h0095FFE3;14'd9743:data <=32'h007CFFD7;
14'd9744:data <=32'h0064FFD2;14'd9745:data <=32'h004FFFD3;14'd9746:data <=32'h003CFFDC;
14'd9747:data <=32'h0032FFE8;14'd9748:data <=32'h0030FFF6;14'd9749:data <=32'h0036FFFF;
14'd9750:data <=32'h00400004;14'd9751:data <=32'h004A0000;14'd9752:data <=32'h0051FFF7;
14'd9753:data <=32'h0053FFEB;14'd9754:data <=32'h004FFFE0;14'd9755:data <=32'h0048FFD9;
14'd9756:data <=32'h003FFFD6;14'd9757:data <=32'h003BFFD8;14'd9758:data <=32'h0038FFDA;
14'd9759:data <=32'h0039FFDB;14'd9760:data <=32'h003DFFD8;14'd9761:data <=32'h0041FFD1;
14'd9762:data <=32'h0041FFC8;14'd9763:data <=32'h003FFFBD;14'd9764:data <=32'h0038FFB3;
14'd9765:data <=32'h002EFFAC;14'd9766:data <=32'h0024FFA7;14'd9767:data <=32'h001AFFA5;
14'd9768:data <=32'h0010FFA6;14'd9769:data <=32'h0007FFA6;14'd9770:data <=32'hFFFFFFA8;
14'd9771:data <=32'hFFF7FFAC;14'd9772:data <=32'hFFEEFFB2;14'd9773:data <=32'hFFEAFFBA;
14'd9774:data <=32'hFFE9FFC4;14'd9775:data <=32'hFFEFFFCE;14'd9776:data <=32'hFFFAFFD3;
14'd9777:data <=32'h0008FFD1;14'd9778:data <=32'h0018FFC6;14'd9779:data <=32'h0024FFB0;
14'd9780:data <=32'h0026FF92;14'd9781:data <=32'h001BFF6F;14'd9782:data <=32'h0002FF4F;
14'd9783:data <=32'hFFDBFF36;14'd9784:data <=32'hFFABFF2A;14'd9785:data <=32'hFF77FF2C;
14'd9786:data <=32'hFF42FF3D;14'd9787:data <=32'hFF13FF5A;14'd9788:data <=32'hFEEAFF83;
14'd9789:data <=32'hFECAFFB6;14'd9790:data <=32'hFEB4FFEF;14'd9791:data <=32'hFEAB0030;
14'd9792:data <=32'hFF280010;14'd9793:data <=32'hFF0A003A;14'd9794:data <=32'hFEF30058;
14'd9795:data <=32'hFED40060;14'd9796:data <=32'hFF1B00C9;14'd9797:data <=32'hFF4C00E6;
14'd9798:data <=32'hFF7A00F4;14'd9799:data <=32'hFFAA00F7;14'd9800:data <=32'hFFD100F0;
14'd9801:data <=32'hFFEF00E6;14'd9802:data <=32'h000900DB;14'd9803:data <=32'h001F00D0;
14'd9804:data <=32'h003500C8;14'd9805:data <=32'h004B00BB;14'd9806:data <=32'h006000AC;
14'd9807:data <=32'h00730099;14'd9808:data <=32'h00820082;14'd9809:data <=32'h008C006A;
14'd9810:data <=32'h00900052;14'd9811:data <=32'h0090003C;14'd9812:data <=32'h00900028;
14'd9813:data <=32'h008C0015;14'd9814:data <=32'h00870001;14'd9815:data <=32'h007EFFED;
14'd9816:data <=32'h0071FFDB;14'd9817:data <=32'h005DFFCC;14'd9818:data <=32'h0044FFC3;
14'd9819:data <=32'h002AFFC3;14'd9820:data <=32'h0012FFCF;14'd9821:data <=32'h0000FFE2;
14'd9822:data <=32'hFFFAFFFB;14'd9823:data <=32'hFFFD0014;14'd9824:data <=32'h000C0028;
14'd9825:data <=32'h00210034;14'd9826:data <=32'h00390037;14'd9827:data <=32'h00500030;
14'd9828:data <=32'h00630024;14'd9829:data <=32'h00700013;14'd9830:data <=32'h0079FFFD;
14'd9831:data <=32'h007CFFE9;14'd9832:data <=32'h007BFFD3;14'd9833:data <=32'h0074FFBF;
14'd9834:data <=32'h0069FFAD;14'd9835:data <=32'h005BFF9E;14'd9836:data <=32'h0048FF93;
14'd9837:data <=32'h0034FF91;14'd9838:data <=32'h0022FF94;14'd9839:data <=32'h0013FF9C;
14'd9840:data <=32'h000EFFA9;14'd9841:data <=32'h000FFFB4;14'd9842:data <=32'h0019FFB9;
14'd9843:data <=32'h0025FFB6;14'd9844:data <=32'h002FFFAA;14'd9845:data <=32'h0034FF94;
14'd9846:data <=32'h002FFF7A;14'd9847:data <=32'h001FFF62;14'd9848:data <=32'h0007FF4D;
14'd9849:data <=32'hFFE8FF41;14'd9850:data <=32'hFFC6FF3C;14'd9851:data <=32'hFFA3FF3F;
14'd9852:data <=32'hFF81FF49;14'd9853:data <=32'hFF63FF59;14'd9854:data <=32'hFF46FF6F;
14'd9855:data <=32'hFF2CFF8A;14'd9856:data <=32'hFF41FF1B;14'd9857:data <=32'hFEF4FF34;
14'd9858:data <=32'hFECCFF62;14'd9859:data <=32'hFF33FFAC;14'd9860:data <=32'hFF58FFFD;
14'd9861:data <=32'hFF61000B;14'd9862:data <=32'hFF690012;14'd9863:data <=32'hFF6D0017;
14'd9864:data <=32'hFF6A001A;14'd9865:data <=32'hFF610022;14'd9866:data <=32'hFF560031;
14'd9867:data <=32'hFF4D004B;14'd9868:data <=32'hFF4B006B;14'd9869:data <=32'hFF540091;
14'd9870:data <=32'hFF6A00B4;14'd9871:data <=32'hFF8900D0;14'd9872:data <=32'hFFB100E5;
14'd9873:data <=32'hFFDA00EF;14'd9874:data <=32'h000600F0;14'd9875:data <=32'h002F00E7;
14'd9876:data <=32'h005600D6;14'd9877:data <=32'h007A00BE;14'd9878:data <=32'h0098009D;
14'd9879:data <=32'h00AD0075;14'd9880:data <=32'h00B60048;14'd9881:data <=32'h00B30019;
14'd9882:data <=32'h009FFFF0;14'd9883:data <=32'h0080FFCF;14'd9884:data <=32'h005BFFBC;
14'd9885:data <=32'h0033FFB8;14'd9886:data <=32'h0011FFC2;14'd9887:data <=32'hFFF6FFD6;
14'd9888:data <=32'hFFE6FFF0;14'd9889:data <=32'hFFE2000B;14'd9890:data <=32'hFFE50024;
14'd9891:data <=32'hFFF00037;14'd9892:data <=32'hFFFF0047;14'd9893:data <=32'h000F0052;
14'd9894:data <=32'h00220058;14'd9895:data <=32'h0035005B;14'd9896:data <=32'h004A005A;
14'd9897:data <=32'h00600054;14'd9898:data <=32'h00750049;14'd9899:data <=32'h00850039;
14'd9900:data <=32'h00930025;14'd9901:data <=32'h009B000F;14'd9902:data <=32'h009FFFFA;
14'd9903:data <=32'h009FFFE6;14'd9904:data <=32'h009EFFD4;14'd9905:data <=32'h009EFFC2;
14'd9906:data <=32'h009DFFAE;14'd9907:data <=32'h009BFF99;14'd9908:data <=32'h0097FF7D;
14'd9909:data <=32'h008AFF60;14'd9910:data <=32'h0074FF42;14'd9911:data <=32'h0054FF2A;
14'd9912:data <=32'h002EFF19;14'd9913:data <=32'h0003FF13;14'd9914:data <=32'hFFD9FF1B;
14'd9915:data <=32'hFFB5FF2C;14'd9916:data <=32'hFF98FF43;14'd9917:data <=32'hFF83FF5E;
14'd9918:data <=32'hFF77FF79;14'd9919:data <=32'hFF6FFF93;14'd9920:data <=32'h001FFEF6;
14'd9921:data <=32'hFFDAFED3;14'd9922:data <=32'hFF8CFEE0;14'd9923:data <=32'hFF6DFFA1;
14'd9924:data <=32'hFF9CFFEE;14'd9925:data <=32'hFFB0FFEF;14'd9926:data <=32'hFFC1FFE5;
14'd9927:data <=32'hFFCBFFD6;14'd9928:data <=32'hFFC9FFC1;14'd9929:data <=32'hFFB8FFAD;
14'd9930:data <=32'hFF9DFFA2;14'd9931:data <=32'hFF7BFFA4;14'd9932:data <=32'hFF58FFB4;
14'd9933:data <=32'hFF3BFFD1;14'd9934:data <=32'hFF29FFF8;14'd9935:data <=32'hFF240022;
14'd9936:data <=32'hFF2A004C;14'd9937:data <=32'hFF3A0074;14'd9938:data <=32'hFF510095;
14'd9939:data <=32'hFF6E00B1;14'd9940:data <=32'hFF9200C5;14'd9941:data <=32'hFFB900D3;
14'd9942:data <=32'hFFE500D8;14'd9943:data <=32'h000F00D0;14'd9944:data <=32'h003600BD;
14'd9945:data <=32'h005400A1;14'd9946:data <=32'h0069007E;14'd9947:data <=32'h00710059;
14'd9948:data <=32'h006D0037;14'd9949:data <=32'h005F001C;14'd9950:data <=32'h004E000A;
14'd9951:data <=32'h003B0000;14'd9952:data <=32'h002BFFFB;14'd9953:data <=32'h001DFFFB;
14'd9954:data <=32'h0012FFFB;14'd9955:data <=32'h0006FFFE;14'd9956:data <=32'hFFFB0001;
14'd9957:data <=32'hFFEE0007;14'd9958:data <=32'hFFE20013;14'd9959:data <=32'hFFD80024;
14'd9960:data <=32'hFFD30039;14'd9961:data <=32'hFFD50052;14'd9962:data <=32'hFFE0006B;
14'd9963:data <=32'hFFF20082;14'd9964:data <=32'h000B0094;14'd9965:data <=32'h002900A1;
14'd9966:data <=32'h004A00A7;14'd9967:data <=32'h006E00A6;14'd9968:data <=32'h0095009E;
14'd9969:data <=32'h00BB008F;14'd9970:data <=32'h00E10074;14'd9971:data <=32'h0104004E;
14'd9972:data <=32'h011F001D;14'd9973:data <=32'h012FFFE2;14'd9974:data <=32'h012DFFA2;
14'd9975:data <=32'h0119FF62;14'd9976:data <=32'h00F3FF2A;14'd9977:data <=32'h00C0FEFF;
14'd9978:data <=32'h0084FEE4;14'd9979:data <=32'h0046FEDD;14'd9980:data <=32'h000EFEE3;
14'd9981:data <=32'hFFDDFEF7;14'd9982:data <=32'hFFB4FF13;14'd9983:data <=32'hFF98FF33;
14'd9984:data <=32'h0053FF61;14'd9985:data <=32'h003EFF3A;14'd9986:data <=32'h000AFF16;
14'd9987:data <=32'hFF8AFF2B;14'd9988:data <=32'hFFA0FF87;14'd9989:data <=32'hFFA5FF9B;
14'd9990:data <=32'hFFAEFFA8;14'd9991:data <=32'hFFB7FFAD;14'd9992:data <=32'hFFBDFFAA;
14'd9993:data <=32'hFFBAFFA1;14'd9994:data <=32'hFFB0FF99;14'd9995:data <=32'hFF9DFF98;
14'd9996:data <=32'hFF89FF9E;14'd9997:data <=32'hFF73FFAE;14'd9998:data <=32'hFF65FFC4;
14'd9999:data <=32'hFF5EFFDD;14'd10000:data <=32'hFF5EFFF6;14'd10001:data <=32'hFF64000B;
14'd10002:data <=32'hFF6C001E;14'd10003:data <=32'hFF76002D;14'd10004:data <=32'hFF7F003A;
14'd10005:data <=32'hFF8A0048;14'd10006:data <=32'hFF970053;14'd10007:data <=32'hFFA7005C;
14'd10008:data <=32'hFFB80062;14'd10009:data <=32'hFFC80061;14'd10010:data <=32'hFFD7005E;
14'd10011:data <=32'hFFE20057;14'd10012:data <=32'hFFE70051;14'd10013:data <=32'hFFEA004E;
14'd10014:data <=32'hFFEC004E;14'd10015:data <=32'hFFF10050;14'd10016:data <=32'hFFFA0052;
14'd10017:data <=32'h00060051;14'd10018:data <=32'h0013004B;14'd10019:data <=32'h001F003F;
14'd10020:data <=32'h0024002D;14'd10021:data <=32'h00210019;14'd10022:data <=32'h00180009;
14'd10023:data <=32'h0004FFFD;14'd10024:data <=32'hFFEDFFFA;14'd10025:data <=32'hFFD40000;
14'd10026:data <=32'hFFC10010;14'd10027:data <=32'hFFB10027;14'd10028:data <=32'hFFA90043;
14'd10029:data <=32'hFFA90063;14'd10030:data <=32'hFFB10084;14'd10031:data <=32'hFFC400A5;
14'd10032:data <=32'hFFDF00C3;14'd10033:data <=32'h000400DC;14'd10034:data <=32'h003300EC;
14'd10035:data <=32'h006800F0;14'd10036:data <=32'h00A200E5;14'd10037:data <=32'h00D800C9;
14'd10038:data <=32'h0106009D;14'd10039:data <=32'h01260064;14'd10040:data <=32'h01360027;
14'd10041:data <=32'h0133FFEA;14'd10042:data <=32'h0122FFB3;14'd10043:data <=32'h0107FF86;
14'd10044:data <=32'h00E6FF64;14'd10045:data <=32'h00C3FF4B;14'd10046:data <=32'h00A0FF39;
14'd10047:data <=32'h007FFF2F;14'd10048:data <=32'h006BFF4E;14'd10049:data <=32'h0057FF38;
14'd10050:data <=32'h004CFF21;14'd10051:data <=32'h007AFF01;14'd10052:data <=32'h0076FF34;
14'd10053:data <=32'h005BFF26;14'd10054:data <=32'h0041FF1D;14'd10055:data <=32'h0023FF16;
14'd10056:data <=32'h0004FF10;14'd10057:data <=32'hFFE2FF0D;14'd10058:data <=32'hFFBAFF11;
14'd10059:data <=32'hFF92FF1F;14'd10060:data <=32'hFF6BFF39;14'd10061:data <=32'hFF4CFF5E;
14'd10062:data <=32'hFF38FF8A;14'd10063:data <=32'hFF33FFBA;14'd10064:data <=32'hFF3CFFE6;
14'd10065:data <=32'hFF4F000A;14'd10066:data <=32'hFF6B0024;14'd10067:data <=32'hFF860032;
14'd10068:data <=32'hFFA10038;14'd10069:data <=32'hFFB80036;14'd10070:data <=32'hFFCA002F;
14'd10071:data <=32'hFFD90027;14'd10072:data <=32'hFFE3001A;14'd10073:data <=32'hFFE8000B;
14'd10074:data <=32'hFFE7FFFD;14'd10075:data <=32'hFFDFFFF0;14'd10076:data <=32'hFFD1FFE8;
14'd10077:data <=32'hFFC0FFE6;14'd10078:data <=32'hFFAEFFED;14'd10079:data <=32'hFFA1FFFC;
14'd10080:data <=32'hFF990011;14'd10081:data <=32'hFF9C0026;14'd10082:data <=32'hFFA80039;
14'd10083:data <=32'hFFB70045;14'd10084:data <=32'hFFC90049;14'd10085:data <=32'hFFDB0045;
14'd10086:data <=32'hFFE5003C;14'd10087:data <=32'hFFE90030;14'd10088:data <=32'hFFE60026;
14'd10089:data <=32'hFFDF001F;14'd10090:data <=32'hFFD50020;14'd10091:data <=32'hFFCB0023;
14'd10092:data <=32'hFFC1002A;14'd10093:data <=32'hFFBB0034;14'd10094:data <=32'hFFB50043;
14'd10095:data <=32'hFFB30054;14'd10096:data <=32'hFFB40067;14'd10097:data <=32'hFFBA007D;
14'd10098:data <=32'hFFC80094;14'd10099:data <=32'hFFDC00AA;14'd10100:data <=32'hFFF700BA;
14'd10101:data <=32'h001900C2;14'd10102:data <=32'h003B00C0;14'd10103:data <=32'h005B00B6;
14'd10104:data <=32'h007600A5;14'd10105:data <=32'h00880091;14'd10106:data <=32'h00960080;
14'd10107:data <=32'h009F0070;14'd10108:data <=32'h00AA0063;14'd10109:data <=32'h00B70057;
14'd10110:data <=32'h00C80049;14'd10111:data <=32'h00DB0035;14'd10112:data <=32'h00F9FFAA;
14'd10113:data <=32'h00EFFF84;14'd10114:data <=32'h00DDFF78;14'd10115:data <=32'h0103FFF8;
14'd10116:data <=32'h0129000B;14'd10117:data <=32'h0132FFD6;14'd10118:data <=32'h0130FF9E;
14'd10119:data <=32'h0120FF66;14'd10120:data <=32'h0106FF2F;14'd10121:data <=32'h00DDFEFD;
14'd10122:data <=32'h00A6FED3;14'd10123:data <=32'h0064FEB8;14'd10124:data <=32'h001BFEAF;
14'd10125:data <=32'hFFD4FEBC;14'd10126:data <=32'hFF94FEDC;14'd10127:data <=32'hFF62FF0C;
14'd10128:data <=32'hFF43FF43;14'd10129:data <=32'hFF37FF7C;14'd10130:data <=32'hFF3AFFB0;
14'd10131:data <=32'hFF48FFDC;14'd10132:data <=32'hFF5EFFFF;14'd10133:data <=32'hFF780018;
14'd10134:data <=32'hFF940028;14'd10135:data <=32'hFFB10030;14'd10136:data <=32'hFFCE0032;
14'd10137:data <=32'hFFE6002B;14'd10138:data <=32'hFFFC001C;14'd10139:data <=32'h00080007;
14'd10140:data <=32'h000CFFF1;14'd10141:data <=32'h0008FFDB;14'd10142:data <=32'hFFFBFFCB;
14'd10143:data <=32'hFFEBFFC1;14'd10144:data <=32'hFFD8FFC0;14'd10145:data <=32'hFFC9FFC3;
14'd10146:data <=32'hFFBFFFCA;14'd10147:data <=32'hFFB7FFD2;14'd10148:data <=32'hFFB3FFD8;
14'd10149:data <=32'hFFAEFFDB;14'd10150:data <=32'hFFA6FFDE;14'd10151:data <=32'hFF9DFFE2;
14'd10152:data <=32'hFF90FFE9;14'd10153:data <=32'hFF84FFF6;14'd10154:data <=32'hFF7A0008;
14'd10155:data <=32'hFF76001D;14'd10156:data <=32'hFF760035;14'd10157:data <=32'hFF7E004B;
14'd10158:data <=32'hFF8A005E;14'd10159:data <=32'hFF98006E;14'd10160:data <=32'hFFAA0078;
14'd10161:data <=32'hFFBB0080;14'd10162:data <=32'hFFCC0085;14'd10163:data <=32'hFFDD0088;
14'd10164:data <=32'hFFEE0087;14'd10165:data <=32'hFFFE0082;14'd10166:data <=32'h000C0079;
14'd10167:data <=32'h0014006D;14'd10168:data <=32'h00160060;14'd10169:data <=32'h00100057;
14'd10170:data <=32'h00050055;14'd10171:data <=32'hFFF9005F;14'd10172:data <=32'hFFF20072;
14'd10173:data <=32'hFFF6008D;14'd10174:data <=32'h000700A8;14'd10175:data <=32'h002400C1;
14'd10176:data <=32'h00B00093;14'd10177:data <=32'h00D00082;14'd10178:data <=32'h00CE006A;
14'd10179:data <=32'h006E009D;14'd10180:data <=32'h00AF00D2;14'd10181:data <=32'h00DB00B8;
14'd10182:data <=32'h01030092;14'd10183:data <=32'h01210064;14'd10184:data <=32'h0136002E;
14'd10185:data <=32'h013FFFF0;14'd10186:data <=32'h0138FFB1;14'd10187:data <=32'h011FFF73;
14'd10188:data <=32'h00F6FF40;14'd10189:data <=32'h00C2FF1B;14'd10190:data <=32'h0088FF07;
14'd10191:data <=32'h0052FF05;14'd10192:data <=32'h0021FF0F;14'd10193:data <=32'hFFFAFF23;
14'd10194:data <=32'hFFDBFF39;14'd10195:data <=32'hFFC6FF52;14'd10196:data <=32'hFFB6FF69;
14'd10197:data <=32'hFFAAFF80;14'd10198:data <=32'hFFA2FF96;14'd10199:data <=32'hFF9DFFAF;
14'd10200:data <=32'hFF9EFFC7;14'd10201:data <=32'hFFA5FFDC;14'd10202:data <=32'hFFB0FFEF;
14'd10203:data <=32'hFFC0FFFB;14'd10204:data <=32'hFFD10002;14'd10205:data <=32'hFFE00004;
14'd10206:data <=32'hFFEC0001;14'd10207:data <=32'hFFF7FFFD;14'd10208:data <=32'h0000FFF8;
14'd10209:data <=32'h0008FFF1;14'd10210:data <=32'h0011FFE8;14'd10211:data <=32'h0019FFDA;
14'd10212:data <=32'h001EFFC7;14'd10213:data <=32'h001CFFB0;14'd10214:data <=32'h0011FF97;
14'd10215:data <=32'hFFFBFF81;14'd10216:data <=32'hFFDDFF6F;14'd10217:data <=32'hFFB7FF6A;
14'd10218:data <=32'hFF8FFF6F;14'd10219:data <=32'hFF6AFF82;14'd10220:data <=32'hFF4CFF9F;
14'd10221:data <=32'hFF37FFC3;14'd10222:data <=32'hFF2DFFEB;14'd10223:data <=32'hFF2D0013;
14'd10224:data <=32'hFF360037;14'd10225:data <=32'hFF460057;14'd10226:data <=32'hFF5D0072;
14'd10227:data <=32'hFF760087;14'd10228:data <=32'hFF930095;14'd10229:data <=32'hFFB2009A;
14'd10230:data <=32'hFFD00095;14'd10231:data <=32'hFFE80089;14'd10232:data <=32'hFFF70077;
14'd10233:data <=32'hFFFC0062;14'd10234:data <=32'hFFF70052;14'd10235:data <=32'hFFE80049;
14'd10236:data <=32'hFFD8004C;14'd10237:data <=32'hFFC8005A;14'd10238:data <=32'hFFC30074;
14'd10239:data <=32'hFFC70091;14'd10240:data <=32'hFFC7008A;14'd10241:data <=32'hFFD500B1;
14'd10242:data <=32'hFFF100BA;14'd10243:data <=32'h001B0086;14'd10244:data <=32'h004600C5;
14'd10245:data <=32'h006300BA;14'd10246:data <=32'h007D00AC;14'd10247:data <=32'h00940098;
14'd10248:data <=32'h00A90081;14'd10249:data <=32'h00BA0066;14'd10250:data <=32'h00C50046;
14'd10251:data <=32'h00C80024;14'd10252:data <=32'h00C20005;14'd10253:data <=32'h00B5FFEB;
14'd10254:data <=32'h00A3FFD7;14'd10255:data <=32'h0093FFCC;14'd10256:data <=32'h0084FFC7;
14'd10257:data <=32'h007DFFC3;14'd10258:data <=32'h007AFFC0;14'd10259:data <=32'h0078FFB5;
14'd10260:data <=32'h0075FFA7;14'd10261:data <=32'h006CFF95;14'd10262:data <=32'h005CFF83;
14'd10263:data <=32'h0047FF77;14'd10264:data <=32'h002EFF6F;14'd10265:data <=32'h0013FF70;
14'd10266:data <=32'hFFFAFF77;14'd10267:data <=32'hFFE6FF83;14'd10268:data <=32'hFFD5FF93;
14'd10269:data <=32'hFFC9FFA6;14'd10270:data <=32'hFFC1FFBA;14'd10271:data <=32'hFFBEFFD0;
14'd10272:data <=32'hFFC3FFE7;14'd10273:data <=32'hFFCEFFFD;14'd10274:data <=32'hFFE1000E;
14'd10275:data <=32'hFFFB0017;14'd10276:data <=32'h00190016;14'd10277:data <=32'h00350009;
14'd10278:data <=32'h004CFFF0;14'd10279:data <=32'h0058FFCE;14'd10280:data <=32'h0057FFA9;
14'd10281:data <=32'h0049FF85;14'd10282:data <=32'h002EFF67;14'd10283:data <=32'h000CFF54;
14'd10284:data <=32'hFFE8FF4B;14'd10285:data <=32'hFFC4FF4C;14'd10286:data <=32'hFFA2FF56;
14'd10287:data <=32'hFF84FF64;14'd10288:data <=32'hFF6CFF79;14'd10289:data <=32'hFF57FF90;
14'd10290:data <=32'hFF46FFAA;14'd10291:data <=32'hFF3BFFC7;14'd10292:data <=32'hFF35FFE5;
14'd10293:data <=32'hFF370003;14'd10294:data <=32'hFF3C001F;14'd10295:data <=32'hFF470035;
14'd10296:data <=32'hFF540046;14'd10297:data <=32'hFF5F0052;14'd10298:data <=32'hFF66005C;
14'd10299:data <=32'hFF6A0069;14'd10300:data <=32'hFF6E0079;14'd10301:data <=32'hFF74008E;
14'd10302:data <=32'hFF7F00A8;14'd10303:data <=32'hFF9400C1;14'd10304:data <=32'hFFA90001;
14'd10305:data <=32'hFF870021;14'd10306:data <=32'hFF7F0052;14'd10307:data <=32'hFFEF00D0;
14'd10308:data <=32'h002A0106;14'd10309:data <=32'h005300ED;14'd10310:data <=32'h007300CD;
14'd10311:data <=32'h008700A9;14'd10312:data <=32'h00930087;14'd10313:data <=32'h00980065;
14'd10314:data <=32'h00960045;14'd10315:data <=32'h008B0028;14'd10316:data <=32'h00790012;
14'd10317:data <=32'h00620002;14'd10318:data <=32'h004B0000;14'd10319:data <=32'h00360008;
14'd10320:data <=32'h002C0018;14'd10321:data <=32'h002C002C;14'd10322:data <=32'h0038003E;
14'd10323:data <=32'h004C0046;14'd10324:data <=32'h00660043;14'd10325:data <=32'h007E0037;
14'd10326:data <=32'h00900020;14'd10327:data <=32'h00990005;14'd10328:data <=32'h0099FFE8;
14'd10329:data <=32'h0091FFCE;14'd10330:data <=32'h0084FFB6;14'd10331:data <=32'h0073FFA4;
14'd10332:data <=32'h005DFF97;14'd10333:data <=32'h0047FF8E;14'd10334:data <=32'h002EFF8B;
14'd10335:data <=32'h0015FF8E;14'd10336:data <=32'hFFFFFF99;14'd10337:data <=32'hFFEEFFAB;
14'd10338:data <=32'hFFE4FFC1;14'd10339:data <=32'hFFE3FFD9;14'd10340:data <=32'hFFEDFFEE;
14'd10341:data <=32'hFFFDFFFC;14'd10342:data <=32'h00110002;14'd10343:data <=32'h0025FFFD;
14'd10344:data <=32'h0036FFF3;14'd10345:data <=32'h0041FFE3;14'd10346:data <=32'h0045FFD2;
14'd10347:data <=32'h0043FFC2;14'd10348:data <=32'h0040FFB4;14'd10349:data <=32'h003CFFA8;
14'd10350:data <=32'h0038FF9C;14'd10351:data <=32'h0033FF8E;14'd10352:data <=32'h002DFF7F;
14'd10353:data <=32'h0021FF6D;14'd10354:data <=32'h0010FF5A;14'd10355:data <=32'hFFF9FF48;
14'd10356:data <=32'hFFDBFF3E;14'd10357:data <=32'hFFBBFF38;14'd10358:data <=32'hFF97FF39;
14'd10359:data <=32'hFF73FF40;14'd10360:data <=32'hFF50FF4D;14'd10361:data <=32'hFF2CFF61;
14'd10362:data <=32'hFF08FF7C;14'd10363:data <=32'hFEE9FFA2;14'd10364:data <=32'hFECCFFCF;
14'd10365:data <=32'hFEBB0008;14'd10366:data <=32'hFEB60049;14'd10367:data <=32'hFEC5008C;
14'd10368:data <=32'hFFAA0003;14'd10369:data <=32'hFF890009;14'd10370:data <=32'hFF5C0025;
14'd10371:data <=32'hFF1000C3;14'd10372:data <=32'hFF580124;14'd10373:data <=32'hFF99012D;
14'd10374:data <=32'hFFD50126;14'd10375:data <=32'h000A0112;14'd10376:data <=32'h003500F8;
14'd10377:data <=32'h005800D8;14'd10378:data <=32'h007000B3;14'd10379:data <=32'h007E008B;
14'd10380:data <=32'h00800064;14'd10381:data <=32'h00760040;14'd10382:data <=32'h00620028;
14'd10383:data <=32'h004A001A;14'd10384:data <=32'h00330018;14'd10385:data <=32'h00220021;
14'd10386:data <=32'h001C002F;14'd10387:data <=32'h001E003E;14'd10388:data <=32'h00280047;
14'd10389:data <=32'h0037004A;14'd10390:data <=32'h00450047;14'd10391:data <=32'h0051003E;
14'd10392:data <=32'h00580033;14'd10393:data <=32'h005B0028;14'd10394:data <=32'h005D001F;
14'd10395:data <=32'h005E0017;14'd10396:data <=32'h0060000F;14'd10397:data <=32'h00600006;
14'd10398:data <=32'h005FFFFC;14'd10399:data <=32'h005CFFF2;14'd10400:data <=32'h0057FFE7;
14'd10401:data <=32'h0050FFE1;14'd10402:data <=32'h0048FFDE;14'd10403:data <=32'h0042FFDD;
14'd10404:data <=32'h003EFFDD;14'd10405:data <=32'h003DFFDD;14'd10406:data <=32'h003DFFDA;
14'd10407:data <=32'h003DFFD6;14'd10408:data <=32'h0039FFD0;14'd10409:data <=32'h0032FFCA;
14'd10410:data <=32'h0029FFC8;14'd10411:data <=32'h001EFFCC;14'd10412:data <=32'h0018FFD4;
14'd10413:data <=32'h0018FFE1;14'd10414:data <=32'h001EFFED;14'd10415:data <=32'h002EFFF6;
14'd10416:data <=32'h0044FFF7;14'd10417:data <=32'h005CFFED;14'd10418:data <=32'h0071FFD8;
14'd10419:data <=32'h0080FFBB;14'd10420:data <=32'h0086FF96;14'd10421:data <=32'h0081FF6F;
14'd10422:data <=32'h0072FF48;14'd10423:data <=32'h0057FF23;14'd10424:data <=32'h0034FF02;
14'd10425:data <=32'h0006FEE8;14'd10426:data <=32'hFFCFFED6;14'd10427:data <=32'hFF90FED2;
14'd10428:data <=32'hFF4DFEDD;14'd10429:data <=32'hFF0CFEFC;14'd10430:data <=32'hFED2FF2E;
14'd10431:data <=32'hFEA7FF70;14'd10432:data <=32'hFF47FF9C;14'd10433:data <=32'hFF1FFFB0;
14'd10434:data <=32'hFEFDFFB9;14'd10435:data <=32'hFEC5FFB4;14'd10436:data <=32'hFEDA002B;
14'd10437:data <=32'hFEF30055;14'd10438:data <=32'hFF0E0077;14'd10439:data <=32'hFF2B008F;
14'd10440:data <=32'hFF4900A4;14'd10441:data <=32'hFF6900B4;14'd10442:data <=32'hFF8A00BE;
14'd10443:data <=32'hFFAA00C2;14'd10444:data <=32'hFFC800BF;14'd10445:data <=32'hFFE300B6;
14'd10446:data <=32'hFFF600AB;14'd10447:data <=32'h000600A0;14'd10448:data <=32'h00110098;
14'd10449:data <=32'h001D0092;14'd10450:data <=32'h002A008D;14'd10451:data <=32'h003B0086;
14'd10452:data <=32'h004D0079;14'd10453:data <=32'h005C0066;14'd10454:data <=32'h0066004E;
14'd10455:data <=32'h00670033;14'd10456:data <=32'h005F001C;14'd10457:data <=32'h004F0009;
14'd10458:data <=32'h003CFFFF;14'd10459:data <=32'h0028FFFD;14'd10460:data <=32'h00190003;
14'd10461:data <=32'h000E000F;14'd10462:data <=32'h0009001B;14'd10463:data <=32'h00090028;
14'd10464:data <=32'h000D0033;14'd10465:data <=32'h0015003E;14'd10466:data <=32'h00210045;
14'd10467:data <=32'h002F004A;14'd10468:data <=32'h0041004C;14'd10469:data <=32'h00530047;
14'd10470:data <=32'h0065003D;14'd10471:data <=32'h0074002C;14'd10472:data <=32'h007D0015;
14'd10473:data <=32'h007EFFFD;14'd10474:data <=32'h0075FFE7;14'd10475:data <=32'h0065FFD7;
14'd10476:data <=32'h0053FFD0;14'd10477:data <=32'h0041FFD1;14'd10478:data <=32'h0036FFDB;
14'd10479:data <=32'h0032FFE8;14'd10480:data <=32'h0038FFF6;14'd10481:data <=32'h0046FFFE;
14'd10482:data <=32'h0058FFFE;14'd10483:data <=32'h006BFFF5;14'd10484:data <=32'h007DFFE6;
14'd10485:data <=32'h0089FFCF;14'd10486:data <=32'h0090FFB5;14'd10487:data <=32'h0093FF99;
14'd10488:data <=32'h008DFF78;14'd10489:data <=32'h0081FF56;14'd10490:data <=32'h006CFF35;
14'd10491:data <=32'h004CFF16;14'd10492:data <=32'h0023FEFE;14'd10493:data <=32'hFFF1FEF1;
14'd10494:data <=32'hFFBDFEF3;14'd10495:data <=32'hFF8BFF02;14'd10496:data <=32'hFFC1FED0;
14'd10497:data <=32'hFF78FEC9;14'd10498:data <=32'hFF49FEDC;14'd10499:data <=32'hFF8DFF2D;
14'd10500:data <=32'hFF89FF7E;14'd10501:data <=32'hFF82FF86;14'd10502:data <=32'hFF77FF8A;
14'd10503:data <=32'hFF68FF8F;14'd10504:data <=32'hFF53FF9A;14'd10505:data <=32'hFF3FFFAB;
14'd10506:data <=32'hFF2DFFC5;14'd10507:data <=32'hFF1FFFE4;14'd10508:data <=32'hFF190006;
14'd10509:data <=32'hFF180028;14'd10510:data <=32'hFF1E004C;14'd10511:data <=32'hFF29006F;
14'd10512:data <=32'hFF3B0093;14'd10513:data <=32'hFF5600B4;14'd10514:data <=32'hFF7900D1;
14'd10515:data <=32'hFFA600E6;14'd10516:data <=32'hFFD900EE;14'd10517:data <=32'h000D00E7;
14'd10518:data <=32'h003D00CF;14'd10519:data <=32'h006200AB;14'd10520:data <=32'h00770080;
14'd10521:data <=32'h007E0053;14'd10522:data <=32'h0076002A;14'd10523:data <=32'h0063000B;
14'd10524:data <=32'h004AFFF5;14'd10525:data <=32'h0030FFE9;14'd10526:data <=32'h0016FFE6;
14'd10527:data <=32'hFFFEFFEA;14'd10528:data <=32'hFFEAFFF5;14'd10529:data <=32'hFFDB0005;
14'd10530:data <=32'hFFCF0018;14'd10531:data <=32'hFFCB002F;14'd10532:data <=32'hFFCF0048;
14'd10533:data <=32'hFFDB005F;14'd10534:data <=32'hFFED0070;14'd10535:data <=32'h0004007D;
14'd10536:data <=32'h001E007F;14'd10537:data <=32'h0036007B;14'd10538:data <=32'h00490072;
14'd10539:data <=32'h00570065;14'd10540:data <=32'h0061005A;14'd10541:data <=32'h00670051;
14'd10542:data <=32'h006F004B;14'd10543:data <=32'h00790046;14'd10544:data <=32'h0086003F;
14'd10545:data <=32'h00970035;14'd10546:data <=32'h00A60024;14'd10547:data <=32'h00B4000C;
14'd10548:data <=32'h00BBFFF0;14'd10549:data <=32'h00BCFFD2;14'd10550:data <=32'h00B5FFB4;
14'd10551:data <=32'h00A9FF99;14'd10552:data <=32'h0099FF84;14'd10553:data <=32'h0085FF70;
14'd10554:data <=32'h0071FF60;14'd10555:data <=32'h0058FF53;14'd10556:data <=32'h003FFF4A;
14'd10557:data <=32'h0022FF46;14'd10558:data <=32'h0007FF4A;14'd10559:data <=32'hFFEEFF57;
14'd10560:data <=32'h00AEFF0F;14'd10561:data <=32'h0082FED6;14'd10562:data <=32'h003DFEC6;
14'd10563:data <=32'hFFEFFF6D;14'd10564:data <=32'hFFFFFFB5;14'd10565:data <=32'h000FFFAD;
14'd10566:data <=32'h0018FF9A;14'd10567:data <=32'h0018FF80;14'd10568:data <=32'h000AFF66;
14'd10569:data <=32'hFFF1FF50;14'd10570:data <=32'hFFCFFF44;14'd10571:data <=32'hFFA9FF41;
14'd10572:data <=32'hFF84FF48;14'd10573:data <=32'hFF5FFF57;14'd10574:data <=32'hFF3DFF70;
14'd10575:data <=32'hFF1EFF91;14'd10576:data <=32'hFF07FFBA;14'd10577:data <=32'hFEF9FFEB;
14'd10578:data <=32'hFEF90020;14'd10579:data <=32'hFF080056;14'd10580:data <=32'hFF260085;
14'd10581:data <=32'hFF4E00A9;14'd10582:data <=32'hFF8100BF;14'd10583:data <=32'hFFB300C3;
14'd10584:data <=32'hFFE100BB;14'd10585:data <=32'h000500A6;14'd10586:data <=32'h001E008C;
14'd10587:data <=32'h002E0071;14'd10588:data <=32'h00350058;14'd10589:data <=32'h00370041;
14'd10590:data <=32'h0035002B;14'd10591:data <=32'h002F0019;14'd10592:data <=32'h00260008;
14'd10593:data <=32'h0018FFFA;14'd10594:data <=32'h0006FFF0;14'd10595:data <=32'hFFF1FFEC;
14'd10596:data <=32'hFFDCFFF0;14'd10597:data <=32'hFFCAFFFA;14'd10598:data <=32'hFFBA0009;
14'd10599:data <=32'hFFB0001C;14'd10600:data <=32'hFFAB0031;14'd10601:data <=32'hFFAA0045;
14'd10602:data <=32'hFFAC005B;14'd10603:data <=32'hFFB10070;14'd10604:data <=32'hFFBA0088;
14'd10605:data <=32'hFFC800A1;14'd10606:data <=32'hFFDE00BB;14'd10607:data <=32'hFFFE00D2;
14'd10608:data <=32'h002700E4;14'd10609:data <=32'h005700EA;14'd10610:data <=32'h008C00E1;
14'd10611:data <=32'h00BF00CA;14'd10612:data <=32'h00EB00A4;14'd10613:data <=32'h010B0072;
14'd10614:data <=32'h011D003D;14'd10615:data <=32'h01200004;14'd10616:data <=32'h0116FFD0;
14'd10617:data <=32'h0101FFA1;14'd10618:data <=32'h00E4FF7A;14'd10619:data <=32'h00C1FF5A;
14'd10620:data <=32'h0099FF44;14'd10621:data <=32'h006FFF38;14'd10622:data <=32'h0043FF38;
14'd10623:data <=32'h001CFF45;14'd10624:data <=32'h00B3FFB5;14'd10625:data <=32'h00B5FF8B;
14'd10626:data <=32'h009BFF59;14'd10627:data <=32'h0017FF4A;14'd10628:data <=32'h0017FF9F;
14'd10629:data <=32'h0020FFA6;14'd10630:data <=32'h002BFFA3;14'd10631:data <=32'h0032FF96;
14'd10632:data <=32'h0031FF86;14'd10633:data <=32'h0028FF75;14'd10634:data <=32'h0016FF66;
14'd10635:data <=32'h0001FF5D;14'd10636:data <=32'hFFEAFF58;14'd10637:data <=32'hFFD4FF59;
14'd10638:data <=32'hFFBCFF5C;14'd10639:data <=32'hFFA4FF63;14'd10640:data <=32'hFF8BFF70;
14'd10641:data <=32'hFF74FF83;14'd10642:data <=32'hFF61FF9C;14'd10643:data <=32'hFF56FFBB;
14'd10644:data <=32'hFF53FFDC;14'd10645:data <=32'hFF59FFFB;14'd10646:data <=32'hFF680013;
14'd10647:data <=32'hFF7A0024;14'd10648:data <=32'hFF8C002D;14'd10649:data <=32'hFF9A0030;
14'd10650:data <=32'hFFA50033;14'd10651:data <=32'hFFAC0035;14'd10652:data <=32'hFFB2003A;
14'd10653:data <=32'hFFBA0041;14'd10654:data <=32'hFFC50047;14'd10655:data <=32'hFFD4004B;
14'd10656:data <=32'hFFE4004B;14'd10657:data <=32'hFFF50043;14'd10658:data <=32'h00020038;
14'd10659:data <=32'h000A0028;14'd10660:data <=32'h000B0016;14'd10661:data <=32'h00060005;
14'd10662:data <=32'hFFFDFFF6;14'd10663:data <=32'hFFEEFFEB;14'd10664:data <=32'hFFDCFFE3;
14'd10665:data <=32'hFFC5FFE0;14'd10666:data <=32'hFFAEFFE3;14'd10667:data <=32'hFF94FFEF;
14'd10668:data <=32'hFF790002;14'd10669:data <=32'hFF630021;14'd10670:data <=32'hFF540049;
14'd10671:data <=32'hFF520079;14'd10672:data <=32'hFF6000AE;14'd10673:data <=32'hFF7E00DE;
14'd10674:data <=32'hFFAC0105;14'd10675:data <=32'hFFE4011E;14'd10676:data <=32'h00220126;
14'd10677:data <=32'h005E011D;14'd10678:data <=32'h00940105;14'd10679:data <=32'h00C100E3;
14'd10680:data <=32'h00E300BB;14'd10681:data <=32'h00FB008D;14'd10682:data <=32'h010A005F;
14'd10683:data <=32'h010F0030;14'd10684:data <=32'h01090003;14'd10685:data <=32'h00FCFFD8;
14'd10686:data <=32'h00E6FFB4;14'd10687:data <=32'h00C9FF99;14'd10688:data <=32'h009CFFBC;
14'd10689:data <=32'h0096FFAE;14'd10690:data <=32'h009DFF9A;14'd10691:data <=32'h00D4FF83;
14'd10692:data <=32'h00C9FFB4;14'd10693:data <=32'h00C4FF9C;14'd10694:data <=32'h00BBFF81;
14'd10695:data <=32'h00ADFF63;14'd10696:data <=32'h0094FF45;14'd10697:data <=32'h0072FF2E;
14'd10698:data <=32'h004AFF20;14'd10699:data <=32'h001FFF20;14'd10700:data <=32'hFFF8FF29;
14'd10701:data <=32'hFFD7FF39;14'd10702:data <=32'hFFBEFF4F;14'd10703:data <=32'hFFAAFF67;
14'd10704:data <=32'hFF9EFF81;14'd10705:data <=32'hFF97FF99;14'd10706:data <=32'hFF95FFB2;
14'd10707:data <=32'hFF98FFCA;14'd10708:data <=32'hFFA2FFDF;14'd10709:data <=32'hFFB1FFEE;
14'd10710:data <=32'hFFC4FFF5;14'd10711:data <=32'hFFD7FFF4;14'd10712:data <=32'hFFE5FFEA;
14'd10713:data <=32'hFFEBFFDB;14'd10714:data <=32'hFFE6FFCC;14'd10715:data <=32'hFFD9FFC0;
14'd10716:data <=32'hFFC8FFBB;14'd10717:data <=32'hFFB5FFC0;14'd10718:data <=32'hFFA5FFCC;
14'd10719:data <=32'hFF9CFFDF;14'd10720:data <=32'hFF9AFFF2;14'd10721:data <=32'hFF9E0003;
14'd10722:data <=32'hFFA90010;14'd10723:data <=32'hFFB50019;14'd10724:data <=32'hFFC2001C;
14'd10725:data <=32'hFFCC001B;14'd10726:data <=32'hFFD50016;14'd10727:data <=32'hFFDC0010;
14'd10728:data <=32'hFFE00007;14'd10729:data <=32'hFFE0FFFB;14'd10730:data <=32'hFFDAFFEE;
14'd10731:data <=32'hFFCDFFE4;14'd10732:data <=32'hFFBAFFDC;14'd10733:data <=32'hFFA2FFDD;
14'd10734:data <=32'hFF88FFE7;14'd10735:data <=32'hFF70FFFD;14'd10736:data <=32'hFF5E001B;
14'd10737:data <=32'hFF58003F;14'd10738:data <=32'hFF5C0065;14'd10739:data <=32'hFF6B0087;
14'd10740:data <=32'hFF8200A3;14'd10741:data <=32'hFF9D00B7;14'd10742:data <=32'hFFBA00C4;
14'd10743:data <=32'hFFD400CC;14'd10744:data <=32'hFFED00D1;14'd10745:data <=32'h000500D3;
14'd10746:data <=32'h001F00D7;14'd10747:data <=32'h003A00D7;14'd10748:data <=32'h005700D3;
14'd10749:data <=32'h007500CA;14'd10750:data <=32'h009000BC;14'd10751:data <=32'h00AA00AA;
14'd10752:data <=32'h00DF0022;14'd10753:data <=32'h00DB0007;14'd10754:data <=32'h00D10007;
14'd10755:data <=32'h00DB0093;14'd10756:data <=32'h00FF00BB;14'd10757:data <=32'h01280090;
14'd10758:data <=32'h01480057;14'd10759:data <=32'h015B0016;14'd10760:data <=32'h015AFFCD;
14'd10761:data <=32'h0146FF87;14'd10762:data <=32'h011EFF4A;14'd10763:data <=32'h00E9FF1B;
14'd10764:data <=32'h00ACFEFF;14'd10765:data <=32'h006EFEF4;14'd10766:data <=32'h0034FEF8;
14'd10767:data <=32'h0001FF08;14'd10768:data <=32'hFFD6FF21;14'd10769:data <=32'hFFB5FF41;
14'd10770:data <=32'hFF9CFF66;14'd10771:data <=32'hFF8FFF8E;14'd10772:data <=32'hFF8DFFB6;
14'd10773:data <=32'hFF98FFDA;14'd10774:data <=32'hFFADFFF8;14'd10775:data <=32'hFFC90009;
14'd10776:data <=32'hFFE7000F;14'd10777:data <=32'h00000006;14'd10778:data <=32'h0014FFF7;
14'd10779:data <=32'h001CFFE2;14'd10780:data <=32'h001BFFCF;14'd10781:data <=32'h0013FFBF;
14'd10782:data <=32'h0007FFB5;14'd10783:data <=32'hFFFAFFB0;14'd10784:data <=32'hFFF1FFB1;
14'd10785:data <=32'hFFE7FFB2;14'd10786:data <=32'hFFE0FFB2;14'd10787:data <=32'hFFDBFFB3;
14'd10788:data <=32'hFFD2FFB3;14'd10789:data <=32'hFFC9FFB2;14'd10790:data <=32'hFFBFFFB6;
14'd10791:data <=32'hFFB6FFBA;14'd10792:data <=32'hFFADFFC1;14'd10793:data <=32'hFFA6FFC9;
14'd10794:data <=32'hFFA0FFD2;14'd10795:data <=32'hFF9BFFD8;14'd10796:data <=32'hFF97FFDF;
14'd10797:data <=32'hFF8FFFE8;14'd10798:data <=32'hFF88FFF1;14'd10799:data <=32'hFF82FFFE;
14'd10800:data <=32'hFF7F0010;14'd10801:data <=32'hFF820022;14'd10802:data <=32'hFF890033;
14'd10803:data <=32'hFF96003F;14'd10804:data <=32'hFFA40045;14'd10805:data <=32'hFFB00043;
14'd10806:data <=32'hFFB7003E;14'd10807:data <=32'hFFB50037;14'd10808:data <=32'hFFAC0033;
14'd10809:data <=32'hFF9E0039;14'd10810:data <=32'hFF900045;14'd10811:data <=32'hFF85005D;
14'd10812:data <=32'hFF80007A;14'd10813:data <=32'hFF85009C;14'd10814:data <=32'hFF9400BD;
14'd10815:data <=32'hFFAB00DF;14'd10816:data <=32'h004B00C7;14'd10817:data <=32'h006100C6;
14'd10818:data <=32'h005C00BB;14'd10819:data <=32'hFFEA00E6;14'd10820:data <=32'h0017013E;
14'd10821:data <=32'h005A0140;14'd10822:data <=32'h009F0130;14'd10823:data <=32'h00DE010F;
14'd10824:data <=32'h011200DB;14'd10825:data <=32'h0135009B;14'd10826:data <=32'h01450055;
14'd10827:data <=32'h01410012;14'd10828:data <=32'h012EFFD8;14'd10829:data <=32'h0110FFA7;
14'd10830:data <=32'h00EEFF81;14'd10831:data <=32'h00C7FF67;14'd10832:data <=32'h009EFF54;
14'd10833:data <=32'h0077FF4A;14'd10834:data <=32'h004FFF48;14'd10835:data <=32'h002AFF4F;
14'd10836:data <=32'h0008FF5E;14'd10837:data <=32'hFFF0FF75;14'd10838:data <=32'hFFE0FF8E;
14'd10839:data <=32'hFFD9FFA7;14'd10840:data <=32'hFFDBFFBD;14'd10841:data <=32'hFFE0FFCD;
14'd10842:data <=32'hFFE9FFD6;14'd10843:data <=32'hFFEFFFDD;14'd10844:data <=32'hFFF4FFE1;
14'd10845:data <=32'hFFF7FFE7;14'd10846:data <=32'hFFFBFFEC;14'd10847:data <=32'h0003FFF2;
14'd10848:data <=32'h000FFFF7;14'd10849:data <=32'h001EFFF7;14'd10850:data <=32'h002FFFF0;
14'd10851:data <=32'h003DFFE1;14'd10852:data <=32'h0046FFCB;14'd10853:data <=32'h0047FFB1;
14'd10854:data <=32'h003FFF97;14'd10855:data <=32'h002FFF7F;14'd10856:data <=32'h0019FF6D;
14'd10857:data <=32'hFFFDFF61;14'd10858:data <=32'hFFE0FF5C;14'd10859:data <=32'hFFC3FF5D;
14'd10860:data <=32'hFFA5FF65;14'd10861:data <=32'hFF89FF73;14'd10862:data <=32'hFF70FF88;
14'd10863:data <=32'hFF5BFFA3;14'd10864:data <=32'hFF4FFFC3;14'd10865:data <=32'hFF4BFFE7;
14'd10866:data <=32'hFF530008;14'd10867:data <=32'hFF650024;14'd10868:data <=32'hFF7E0037;
14'd10869:data <=32'hFF99003D;14'd10870:data <=32'hFFAF0037;14'd10871:data <=32'hFFBE0029;
14'd10872:data <=32'hFFC20017;14'd10873:data <=32'hFFBA0008;14'd10874:data <=32'hFFA90000;
14'd10875:data <=32'hFF930000;14'd10876:data <=32'hFF7E000B;14'd10877:data <=32'hFF6B001E;
14'd10878:data <=32'hFF5D0039;14'd10879:data <=32'hFF570058;14'd10880:data <=32'hFF740059;
14'd10881:data <=32'hFF66007D;14'd10882:data <=32'hFF6D0090;14'd10883:data <=32'hFF8A0072;
14'd10884:data <=32'hFF9600D3;14'd10885:data <=32'hFFBA00E8;14'd10886:data <=32'hFFE400F6;
14'd10887:data <=32'h001100F8;14'd10888:data <=32'h003C00EC;14'd10889:data <=32'h006000D6;
14'd10890:data <=32'h007C00BA;14'd10891:data <=32'h008D009C;14'd10892:data <=32'h00940081;
14'd10893:data <=32'h0098006B;14'd10894:data <=32'h009A0059;14'd10895:data <=32'h009E0049;
14'd10896:data <=32'h00A30039;14'd10897:data <=32'h00A80025;14'd10898:data <=32'h00AA0010;
14'd10899:data <=32'h00A6FFFA;14'd10900:data <=32'h00A1FFE3;14'd10901:data <=32'h0096FFD1;
14'd10902:data <=32'h0089FFC0;14'd10903:data <=32'h007BFFB3;14'd10904:data <=32'h006DFFA6;
14'd10905:data <=32'h005BFF9B;14'd10906:data <=32'h0047FF93;14'd10907:data <=32'h0030FF8D;
14'd10908:data <=32'h0017FF8E;14'd10909:data <=32'hFFFDFF97;14'd10910:data <=32'hFFE7FFAB;
14'd10911:data <=32'hFFD8FFC5;14'd10912:data <=32'hFFD4FFE3;14'd10913:data <=32'hFFDE0001;
14'd10914:data <=32'hFFF1001A;14'd10915:data <=32'h000E0028;14'd10916:data <=32'h002C0029;
14'd10917:data <=32'h004B0020;14'd10918:data <=32'h0064000C;14'd10919:data <=32'h0075FFF1;
14'd10920:data <=32'h007EFFD2;14'd10921:data <=32'h007EFFB2;14'd10922:data <=32'h0076FF93;
14'd10923:data <=32'h0066FF76;14'd10924:data <=32'h004FFF5C;14'd10925:data <=32'h0034FF48;
14'd10926:data <=32'h0012FF3B;14'd10927:data <=32'hFFEEFF35;14'd10928:data <=32'hFFC9FF3B;
14'd10929:data <=32'hFFA8FF49;14'd10930:data <=32'hFF8DFF60;14'd10931:data <=32'hFF7CFF79;
14'd10932:data <=32'hFF73FF93;14'd10933:data <=32'hFF72FFA9;14'd10934:data <=32'hFF74FFB7;
14'd10935:data <=32'hFF75FFC1;14'd10936:data <=32'hFF73FFC7;14'd10937:data <=32'hFF6BFFCB;
14'd10938:data <=32'hFF5FFFD4;14'd10939:data <=32'hFF52FFE3;14'd10940:data <=32'hFF46FFF7;
14'd10941:data <=32'hFF400011;14'd10942:data <=32'hFF3F002B;14'd10943:data <=32'hFF440047;
14'd10944:data <=32'hFF9FFFA9;14'd10945:data <=32'hFF67FFAF;14'd10946:data <=32'hFF40FFD5;
14'd10947:data <=32'hFF74006C;14'd10948:data <=32'hFF8400C0;14'd10949:data <=32'hFFAA00C9;
14'd10950:data <=32'hFFD000CA;14'd10951:data <=32'hFFF200C1;14'd10952:data <=32'h001100AE;
14'd10953:data <=32'h00270094;14'd10954:data <=32'h00310077;14'd10955:data <=32'h002E005D;
14'd10956:data <=32'h0022004C;14'd10957:data <=32'h00130046;14'd10958:data <=32'h0004004B;
14'd10959:data <=32'hFFFD0057;14'd10960:data <=32'hFFFF0069;14'd10961:data <=32'h000B0078;
14'd10962:data <=32'h001C0083;14'd10963:data <=32'h00330088;14'd10964:data <=32'h004B0085;
14'd10965:data <=32'h0062007D;14'd10966:data <=32'h00780070;14'd10967:data <=32'h008D005E;
14'd10968:data <=32'h009D0045;14'd10969:data <=32'h00A80029;14'd10970:data <=32'h00AB0007;
14'd10971:data <=32'h00A4FFE5;14'd10972:data <=32'h0092FFC6;14'd10973:data <=32'h0078FFAE;
14'd10974:data <=32'h0057FFA0;14'd10975:data <=32'h0034FF9F;14'd10976:data <=32'h0017FFAA;
14'd10977:data <=32'h0000FFBE;14'd10978:data <=32'hFFF5FFD7;14'd10979:data <=32'hFFF3FFF0;
14'd10980:data <=32'hFFFC0004;14'd10981:data <=32'h00090014;14'd10982:data <=32'h0019001B;
14'd10983:data <=32'h002B001F;14'd10984:data <=32'h003B001E;14'd10985:data <=32'h004A001A;
14'd10986:data <=32'h00590012;14'd10987:data <=32'h00690007;14'd10988:data <=32'h0076FFF7;
14'd10989:data <=32'h0082FFE4;14'd10990:data <=32'h0088FFCD;14'd10991:data <=32'h008AFFB3;
14'd10992:data <=32'h0084FF99;14'd10993:data <=32'h0079FF81;14'd10994:data <=32'h006BFF6A;
14'd10995:data <=32'h005BFF58;14'd10996:data <=32'h0049FF45;14'd10997:data <=32'h0035FF34;
14'd10998:data <=32'h001DFF21;14'd10999:data <=32'h0000FF0F;14'd11000:data <=32'hFFD9FF00;
14'd11001:data <=32'hFFABFEF9;14'd11002:data <=32'hFF77FEFF;14'd11003:data <=32'hFF41FF12;
14'd11004:data <=32'hFF11FF36;14'd11005:data <=32'hFEE9FF66;14'd11006:data <=32'hFED1FF9F;
14'd11007:data <=32'hFEC7FFDA;14'd11008:data <=32'hFFD9FFAC;14'd11009:data <=32'hFFB2FF93;
14'd11010:data <=32'hFF73FF8D;14'd11011:data <=32'hFEE50010;14'd11012:data <=32'hFEF20084;
14'd11013:data <=32'hFF1D00AB;14'd11014:data <=32'hFF5000C5;14'd11015:data <=32'hFF8300D3;
14'd11016:data <=32'hFFB700CE;14'd11017:data <=32'hFFE500BC;14'd11018:data <=32'h0005009E;
14'd11019:data <=32'h0016007B;14'd11020:data <=32'h0019005C;14'd11021:data <=32'h000F0044;
14'd11022:data <=32'hFFFE0036;14'd11023:data <=32'hFFED0034;14'd11024:data <=32'hFFE2003B;
14'd11025:data <=32'hFFDB0046;14'd11026:data <=32'hFFDC0053;14'd11027:data <=32'hFFE20060;
14'd11028:data <=32'hFFEA006A;14'd11029:data <=32'hFFF50071;14'd11030:data <=32'h00040077;
14'd11031:data <=32'h0014007B;14'd11032:data <=32'h0026007C;14'd11033:data <=32'h003A0078;
14'd11034:data <=32'h004D006E;14'd11035:data <=32'h005E005E;14'd11036:data <=32'h00680049;
14'd11037:data <=32'h006A0032;14'd11038:data <=32'h0065001F;14'd11039:data <=32'h005C0010;
14'd11040:data <=32'h00500006;14'd11041:data <=32'h00460004;14'd11042:data <=32'h00410005;
14'd11043:data <=32'h003E0006;14'd11044:data <=32'h003E0006;14'd11045:data <=32'h003D0003;
14'd11046:data <=32'h003BFFFE;14'd11047:data <=32'h0038FFF9;14'd11048:data <=32'h0030FFF7;
14'd11049:data <=32'h0026FFF8;14'd11050:data <=32'h001F0000;14'd11051:data <=32'h001C000B;
14'd11052:data <=32'h001F001A;14'd11053:data <=32'h00280027;14'd11054:data <=32'h00380031;
14'd11055:data <=32'h004C0037;14'd11056:data <=32'h00620036;14'd11057:data <=32'h007C0031;
14'd11058:data <=32'h00960023;14'd11059:data <=32'h00AF0010;14'd11060:data <=32'h00C6FFF4;
14'd11061:data <=32'h00DAFFCE;14'd11062:data <=32'h00E6FF9F;14'd11063:data <=32'h00E6FF68;
14'd11064:data <=32'h00D7FF2C;14'd11065:data <=32'h00B4FEF3;14'd11066:data <=32'h007FFEC2;
14'd11067:data <=32'h003BFEA1;14'd11068:data <=32'hFFF1FE94;14'd11069:data <=32'hFFA4FE9A;
14'd11070:data <=32'hFF5DFEB6;14'd11071:data <=32'hFF22FEE1;14'd11072:data <=32'hFFBAFF5C;
14'd11073:data <=32'hFF98FF4B;14'd11074:data <=32'hFF74FF30;14'd11075:data <=32'hFF21FF0A;
14'd11076:data <=32'hFEF8FF7D;14'd11077:data <=32'hFEF1FFB0;14'd11078:data <=32'hFEF6FFDF;
14'd11079:data <=32'hFF04000C;14'd11080:data <=32'hFF1C002F;14'd11081:data <=32'hFF380048;
14'd11082:data <=32'hFF550056;14'd11083:data <=32'hFF6D005C;14'd11084:data <=32'hFF7F005D;
14'd11085:data <=32'hFF8B005E;14'd11086:data <=32'hFF930062;14'd11087:data <=32'hFF9B006B;
14'd11088:data <=32'hFFA60075;14'd11089:data <=32'hFFB8007E;14'd11090:data <=32'hFFCC0084;
14'd11091:data <=32'hFFE20082;14'd11092:data <=32'hFFF6007C;14'd11093:data <=32'h0005006F;
14'd11094:data <=32'h000F0063;14'd11095:data <=32'h00140056;14'd11096:data <=32'h0017004A;
14'd11097:data <=32'h00160041;14'd11098:data <=32'h00150039;14'd11099:data <=32'h00130032;
14'd11100:data <=32'h000D002C;14'd11101:data <=32'h00080029;14'd11102:data <=32'hFFFF0029;
14'd11103:data <=32'hFFF7002E;14'd11104:data <=32'hFFF10039;14'd11105:data <=32'hFFF10047;
14'd11106:data <=32'hFFF90055;14'd11107:data <=32'h00060063;14'd11108:data <=32'h001B0068;
14'd11109:data <=32'h00310066;14'd11110:data <=32'h0045005B;14'd11111:data <=32'h0052004A;
14'd11112:data <=32'h00580035;14'd11113:data <=32'h00550023;14'd11114:data <=32'h004B0016;
14'd11115:data <=32'h003F000E;14'd11116:data <=32'h0032000F;14'd11117:data <=32'h00280015;
14'd11118:data <=32'h00230020;14'd11119:data <=32'h0023002C;14'd11120:data <=32'h002A003A;
14'd11121:data <=32'h00350046;14'd11122:data <=32'h00460050;14'd11123:data <=32'h005D0057;
14'd11124:data <=32'h00790059;14'd11125:data <=32'h009B0050;14'd11126:data <=32'h00BD003E;
14'd11127:data <=32'h00DD001E;14'd11128:data <=32'h00F5FFF3;14'd11129:data <=32'h00FFFFBE;
14'd11130:data <=32'h00F9FF85;14'd11131:data <=32'h00E4FF4F;14'd11132:data <=32'h00C0FF22;
14'd11133:data <=32'h0093FF01;14'd11134:data <=32'h0061FEEE;14'd11135:data <=32'h0031FEE7;
14'd11136:data <=32'h0063FEEB;14'd11137:data <=32'h0034FEC1;14'd11138:data <=32'h000FFEB0;
14'd11139:data <=32'h002FFEF0;14'd11140:data <=32'hFFFDFF2D;14'd11141:data <=32'hFFE5FF2C;
14'd11142:data <=32'hFFCBFF2F;14'd11143:data <=32'hFFB1FF35;14'd11144:data <=32'hFF9AFF3F;
14'd11145:data <=32'hFF83FF4A;14'd11146:data <=32'hFF6CFF56;14'd11147:data <=32'hFF55FF66;
14'd11148:data <=32'hFF3CFF7A;14'd11149:data <=32'hFF22FF93;14'd11150:data <=32'hFF0DFFB7;
14'd11151:data <=32'hFEFEFFE4;14'd11152:data <=32'hFEFD0017;14'd11153:data <=32'hFF0A004B;
14'd11154:data <=32'hFF250077;14'd11155:data <=32'hFF4D009B;14'd11156:data <=32'hFF7B00AF;
14'd11157:data <=32'hFFAA00B6;14'd11158:data <=32'hFFD600AF;14'd11159:data <=32'hFFFA009F;
14'd11160:data <=32'h00150089;14'd11161:data <=32'h0029006E;14'd11162:data <=32'h00350052;
14'd11163:data <=32'h00390035;14'd11164:data <=32'h00330019;14'd11165:data <=32'h00260000;
14'd11166:data <=32'h0010FFEE;14'd11167:data <=32'hFFF7FFE4;14'd11168:data <=32'hFFDAFFE6;
14'd11169:data <=32'hFFC0FFF3;14'd11170:data <=32'hFFAF0008;14'd11171:data <=32'hFFA60023;
14'd11172:data <=32'hFFA8003E;14'd11173:data <=32'hFFB30055;14'd11174:data <=32'hFFC50067;
14'd11175:data <=32'hFFD6006F;14'd11176:data <=32'hFFE80073;14'd11177:data <=32'hFFF60071;
14'd11178:data <=32'hFFFF0071;14'd11179:data <=32'h00090070;14'd11180:data <=32'h00100072;
14'd11181:data <=32'h00190075;14'd11182:data <=32'h00240078;14'd11183:data <=32'h0032007A;
14'd11184:data <=32'h00410079;14'd11185:data <=32'h00510075;14'd11186:data <=32'h0060006F;
14'd11187:data <=32'h006D0068;14'd11188:data <=32'h007D0060;14'd11189:data <=32'h008C0057;
14'd11190:data <=32'h009D0049;14'd11191:data <=32'h00AD0036;14'd11192:data <=32'h00BB001D;
14'd11193:data <=32'h00C2FFFF;14'd11194:data <=32'h00C2FFE0;14'd11195:data <=32'h00B6FFC1;
14'd11196:data <=32'h00A5FFA9;14'd11197:data <=32'h008EFF99;14'd11198:data <=32'h0078FF91;
14'd11199:data <=32'h0069FF92;14'd11200:data <=32'h011EFF8E;14'd11201:data <=32'h0119FF48;
14'd11202:data <=32'h00F2FF1B;14'd11203:data <=32'h007EFF91;14'd11204:data <=32'h006EFFC7;
14'd11205:data <=32'h007AFFB6;14'd11206:data <=32'h0080FFA0;14'd11207:data <=32'h0080FF82;
14'd11208:data <=32'h0079FF66;14'd11209:data <=32'h006AFF47;14'd11210:data <=32'h0053FF29;
14'd11211:data <=32'h0034FF0D;14'd11212:data <=32'h0009FEF8;14'd11213:data <=32'hFFD4FEEE;
14'd11214:data <=32'hFF99FEF3;14'd11215:data <=32'hFF60FF08;14'd11216:data <=32'hFF2FFF2F;
14'd11217:data <=32'hFF0AFF64;14'd11218:data <=32'hFEF7FF9E;14'd11219:data <=32'hFEF7FFDB;
14'd11220:data <=32'hFF060010;14'd11221:data <=32'hFF20003D;14'd11222:data <=32'hFF42005D;
14'd11223:data <=32'hFF670073;14'd11224:data <=32'hFF8C007F;14'd11225:data <=32'hFFAF0082;
14'd11226:data <=32'hFFD1007F;14'd11227:data <=32'hFFF00074;14'd11228:data <=32'h00090061;
14'd11229:data <=32'h001B0049;14'd11230:data <=32'h0024002D;14'd11231:data <=32'h00230010;
14'd11232:data <=32'h0019FFF8;14'd11233:data <=32'h0008FFE6;14'd11234:data <=32'hFFF4FFDD;
14'd11235:data <=32'hFFE0FFDA;14'd11236:data <=32'hFFCDFFDE;14'd11237:data <=32'hFFBFFFE3;
14'd11238:data <=32'hFFB2FFEB;14'd11239:data <=32'hFFA6FFF3;14'd11240:data <=32'hFF9AFFFD;
14'd11241:data <=32'hFF8D0008;14'd11242:data <=32'hFF7E001B;14'd11243:data <=32'hFF720034;
14'd11244:data <=32'hFF6C0053;14'd11245:data <=32'hFF6E0077;14'd11246:data <=32'hFF7C009C;
14'd11247:data <=32'hFF9300BE;14'd11248:data <=32'hFFB700DB;14'd11249:data <=32'hFFDF00ED;
14'd11250:data <=32'h000B00F5;14'd11251:data <=32'h003600F4;14'd11252:data <=32'h006200E8;
14'd11253:data <=32'h008900D6;14'd11254:data <=32'h00AD00BB;14'd11255:data <=32'h00CB0098;
14'd11256:data <=32'h00E00070;14'd11257:data <=32'h00EC0041;14'd11258:data <=32'h00E90012;
14'd11259:data <=32'h00DAFFE7;14'd11260:data <=32'h00BFFFC4;14'd11261:data <=32'h009CFFAE;
14'd11262:data <=32'h0078FFA8;14'd11263:data <=32'h005AFFAF;14'd11264:data <=32'h00C50045;
14'd11265:data <=32'h00E70029;14'd11266:data <=32'h00F0FFF1;14'd11267:data <=32'h007AFFB1;
14'd11268:data <=32'h0062FFF4;14'd11269:data <=32'h006EFFF3;14'd11270:data <=32'h007AFFEB;
14'd11271:data <=32'h0086FFDE;14'd11272:data <=32'h008EFFCC;14'd11273:data <=32'h0094FFB8;
14'd11274:data <=32'h0096FF9E;14'd11275:data <=32'h0091FF7F;14'd11276:data <=32'h0083FF60;
14'd11277:data <=32'h006BFF41;14'd11278:data <=32'h0047FF2A;14'd11279:data <=32'h001EFF1E;
14'd11280:data <=32'hFFF0FF1D;14'd11281:data <=32'hFFC7FF2C;14'd11282:data <=32'hFFA5FF43;
14'd11283:data <=32'hFF8EFF60;14'd11284:data <=32'hFF80FF7D;14'd11285:data <=32'hFF79FF99;
14'd11286:data <=32'hFF79FFB1;14'd11287:data <=32'hFF7BFFC4;14'd11288:data <=32'hFF7CFFD7;
14'd11289:data <=32'hFF7FFFE8;14'd11290:data <=32'hFF85FFFA;14'd11291:data <=32'hFF8E000C;
14'd11292:data <=32'hFF9B001B;14'd11293:data <=32'hFFAA0024;14'd11294:data <=32'hFFBB002B;
14'd11295:data <=32'hFFCC002A;14'd11296:data <=32'hFFDB0028;14'd11297:data <=32'hFFE70021;
14'd11298:data <=32'hFFF00019;14'd11299:data <=32'hFFF80011;14'd11300:data <=32'hFFFE0007;
14'd11301:data <=32'h0005FFF8;14'd11302:data <=32'h0006FFE5;14'd11303:data <=32'h0001FFD1;
14'd11304:data <=32'hFFF4FFBB;14'd11305:data <=32'hFFDCFFA6;14'd11306:data <=32'hFFBBFF9B;
14'd11307:data <=32'hFF94FF9B;14'd11308:data <=32'hFF69FFA8;14'd11309:data <=32'hFF43FFC5;
14'd11310:data <=32'hFF25FFEE;14'd11311:data <=32'hFF15001F;14'd11312:data <=32'hFF120055;
14'd11313:data <=32'hFF1F008A;14'd11314:data <=32'hFF3700B9;14'd11315:data <=32'hFF5B00E2;
14'd11316:data <=32'hFF860101;14'd11317:data <=32'hFFB70117;14'd11318:data <=32'hFFEB0123;
14'd11319:data <=32'h00200120;14'd11320:data <=32'h00550112;14'd11321:data <=32'h008400F6;
14'd11322:data <=32'h00AB00D1;14'd11323:data <=32'h00C200A5;14'd11324:data <=32'h00CC0077;
14'd11325:data <=32'h00C8004D;14'd11326:data <=32'h00BA002D;14'd11327:data <=32'h00A80019;
14'd11328:data <=32'h00700033;14'd11329:data <=32'h00790036;14'd11330:data <=32'h00960031;
14'd11331:data <=32'h00DB001C;14'd11332:data <=32'h00C50042;14'd11333:data <=32'h00CF0027;
14'd11334:data <=32'h00D50009;14'd11335:data <=32'h00D3FFEA;14'd11336:data <=32'h00CBFFCC;
14'd11337:data <=32'h00BDFFB3;14'd11338:data <=32'h00ADFF9C;14'd11339:data <=32'h009AFF88;
14'd11340:data <=32'h0085FF76;14'd11341:data <=32'h006BFF69;14'd11342:data <=32'h004FFF60;
14'd11343:data <=32'h0030FF5D;14'd11344:data <=32'h0012FF65;14'd11345:data <=32'hFFF9FF75;
14'd11346:data <=32'hFFE9FF8B;14'd11347:data <=32'hFFE4FFA1;14'd11348:data <=32'hFFE7FFB5;
14'd11349:data <=32'hFFF1FFC1;14'd11350:data <=32'hFFFCFFC4;14'd11351:data <=32'h0005FFBE;
14'd11352:data <=32'h0007FFB4;14'd11353:data <=32'h0002FFAA;14'd11354:data <=32'hFFF7FFA2;
14'd11355:data <=32'hFFEAFF9F;14'd11356:data <=32'hFFDCFFA0;14'd11357:data <=32'hFFCFFFA7;
14'd11358:data <=32'hFFC3FFB0;14'd11359:data <=32'hFFBBFFBA;14'd11360:data <=32'hFFB5FFC7;
14'd11361:data <=32'hFFB1FFD4;14'd11362:data <=32'hFFB1FFE4;14'd11363:data <=32'hFFB7FFF3;
14'd11364:data <=32'hFFC20000;14'd11365:data <=32'hFFD20009;14'd11366:data <=32'hFFE50009;
14'd11367:data <=32'hFFF80001;14'd11368:data <=32'h0007FFEF;14'd11369:data <=32'h000CFFD7;
14'd11370:data <=32'h0007FFBB;14'd11371:data <=32'hFFF5FFA2;14'd11372:data <=32'hFFDAFF90;
14'd11373:data <=32'hFFB8FF89;14'd11374:data <=32'hFF94FF8D;14'd11375:data <=32'hFF74FF9C;
14'd11376:data <=32'hFF59FFB3;14'd11377:data <=32'hFF44FFCF;14'd11378:data <=32'hFF37FFEF;
14'd11379:data <=32'hFF30000F;14'd11380:data <=32'hFF2F0031;14'd11381:data <=32'hFF320052;
14'd11382:data <=32'hFF3C0074;14'd11383:data <=32'hFF4D0094;14'd11384:data <=32'hFF6400B0;
14'd11385:data <=32'hFF8000C7;14'd11386:data <=32'hFFA100D6;14'd11387:data <=32'hFFBF00DE;
14'd11388:data <=32'hFFDB00E0;14'd11389:data <=32'hFFF400E0;14'd11390:data <=32'h000A00E0;
14'd11391:data <=32'h002000E3;14'd11392:data <=32'h007B006E;14'd11393:data <=32'h007B0066;
14'd11394:data <=32'h00750073;14'd11395:data <=32'h00680101;14'd11396:data <=32'h00810132;
14'd11397:data <=32'h00BC0116;14'd11398:data <=32'h00F100ED;14'd11399:data <=32'h011700B6;
14'd11400:data <=32'h012D0079;14'd11401:data <=32'h0135003C;14'd11402:data <=32'h012F0002;
14'd11403:data <=32'h011DFFCD;14'd11404:data <=32'h0101FF9C;14'd11405:data <=32'h00DDFF74;
14'd11406:data <=32'h00AFFF57;14'd11407:data <=32'h007EFF47;14'd11408:data <=32'h004BFF45;
14'd11409:data <=32'h001BFF53;14'd11410:data <=32'hFFF6FF6E;14'd11411:data <=32'hFFDFFF91;
14'd11412:data <=32'hFFD8FFB6;14'd11413:data <=32'hFFDDFFD6;14'd11414:data <=32'hFFEEFFED;
14'd11415:data <=32'h0004FFF8;14'd11416:data <=32'h0017FFFA;14'd11417:data <=32'h0028FFF3;
14'd11418:data <=32'h0031FFE8;14'd11419:data <=32'h0037FFDC;14'd11420:data <=32'h0037FFCF;
14'd11421:data <=32'h0035FFC4;14'd11422:data <=32'h0030FFB9;14'd11423:data <=32'h0029FFB0;
14'd11424:data <=32'h0020FFA7;14'd11425:data <=32'h0015FFA2;14'd11426:data <=32'h0007FF9F;
14'd11427:data <=32'hFFFAFFA0;14'd11428:data <=32'hFFEEFFA6;14'd11429:data <=32'hFFE7FFAD;
14'd11430:data <=32'hFFE4FFB6;14'd11431:data <=32'hFFE6FFBB;14'd11432:data <=32'hFFE8FFBC;
14'd11433:data <=32'hFFEAFFB9;14'd11434:data <=32'hFFE9FFB2;14'd11435:data <=32'hFFE2FFAB;
14'd11436:data <=32'hFFD6FFA4;14'd11437:data <=32'hFFC7FFA4;14'd11438:data <=32'hFFB8FFA9;
14'd11439:data <=32'hFFACFFB3;14'd11440:data <=32'hFFA5FFBE;14'd11441:data <=32'hFFA3FFC9;
14'd11442:data <=32'hFFA2FFD1;14'd11443:data <=32'hFFA5FFD4;14'd11444:data <=32'hFFA2FFD4;
14'd11445:data <=32'hFF9CFFD2;14'd11446:data <=32'hFF92FFD0;14'd11447:data <=32'hFF83FFD2;
14'd11448:data <=32'hFF72FFD9;14'd11449:data <=32'hFF62FFE4;14'd11450:data <=32'hFF51FFF4;
14'd11451:data <=32'hFF420007;14'd11452:data <=32'hFF33001F;14'd11453:data <=32'hFF25003F;
14'd11454:data <=32'hFF1C0065;14'd11455:data <=32'hFF1A0094;14'd11456:data <=32'hFFD000B3;
14'd11457:data <=32'hFFD900C0;14'd11458:data <=32'hFFD000C0;14'd11459:data <=32'hFF5200DB;
14'd11460:data <=32'hFF640142;14'd11461:data <=32'hFFA9015F;14'd11462:data <=32'hFFF30169;
14'd11463:data <=32'h003D015F;14'd11464:data <=32'h007B0145;14'd11465:data <=32'h00B1011F;
14'd11466:data <=32'h00DB00F0;14'd11467:data <=32'h00FA00BD;14'd11468:data <=32'h010C0085;
14'd11469:data <=32'h0112004C;14'd11470:data <=32'h010B0014;14'd11471:data <=32'h00F6FFE2;
14'd11472:data <=32'h00D7FFBA;14'd11473:data <=32'h00AFFF9F;14'd11474:data <=32'h0086FF92;
14'd11475:data <=32'h0060FF92;14'd11476:data <=32'h0041FF9C;14'd11477:data <=32'h002CFFAA;
14'd11478:data <=32'h0021FFB9;14'd11479:data <=32'h001CFFC5;14'd11480:data <=32'h0019FFCE;
14'd11481:data <=32'h0017FFD5;14'd11482:data <=32'h0014FFDA;14'd11483:data <=32'h0011FFE1;
14'd11484:data <=32'h000FFFEA;14'd11485:data <=32'h0011FFF4;14'd11486:data <=32'h0018FFFD;
14'd11487:data <=32'h00230004;14'd11488:data <=32'h002F0004;14'd11489:data <=32'h003D0001;
14'd11490:data <=32'h0048FFF9;14'd11491:data <=32'h0052FFED;14'd11492:data <=32'h0058FFE0;
14'd11493:data <=32'h005BFFD0;14'd11494:data <=32'h005DFFC0;14'd11495:data <=32'h005CFFAF;
14'd11496:data <=32'h0056FF9C;14'd11497:data <=32'h004DFF86;14'd11498:data <=32'h003CFF72;
14'd11499:data <=32'h0025FF62;14'd11500:data <=32'h0006FF59;14'd11501:data <=32'hFFE5FF57;
14'd11502:data <=32'hFFC6FF61;14'd11503:data <=32'hFFADFF76;14'd11504:data <=32'hFF9CFF90;
14'd11505:data <=32'hFF95FFAC;14'd11506:data <=32'hFF9BFFC4;14'd11507:data <=32'hFFA7FFD6;
14'd11508:data <=32'hFFB6FFDD;14'd11509:data <=32'hFFC5FFDC;14'd11510:data <=32'hFFCEFFD5;
14'd11511:data <=32'hFFD2FFC7;14'd11512:data <=32'hFFCFFFBB;14'd11513:data <=32'hFFC5FFAD;
14'd11514:data <=32'hFFB5FFA0;14'd11515:data <=32'hFF9FFF98;14'd11516:data <=32'hFF83FF94;
14'd11517:data <=32'hFF61FF97;14'd11518:data <=32'hFF3BFFA6;14'd11519:data <=32'hFF15FFC2;
14'd11520:data <=32'hFF43FFED;14'd11521:data <=32'hFF1F000C;14'd11522:data <=32'hFF130023;
14'd11523:data <=32'hFF270011;14'd11524:data <=32'hFF0C0078;14'd11525:data <=32'hFF2800A4;
14'd11526:data <=32'hFF4C00C6;14'd11527:data <=32'hFF7400DA;14'd11528:data <=32'hFF9C00E6;
14'd11529:data <=32'hFFC000E9;14'd11530:data <=32'hFFE100E8;14'd11531:data <=32'h000200E3;
14'd11532:data <=32'h001F00DC;14'd11533:data <=32'h003D00CF;14'd11534:data <=32'h005600BD;
14'd11535:data <=32'h006B00A7;14'd11536:data <=32'h007A008F;14'd11537:data <=32'h00820078;
14'd11538:data <=32'h00870062;14'd11539:data <=32'h00890051;14'd11540:data <=32'h008B0041;
14'd11541:data <=32'h008E0032;14'd11542:data <=32'h00930020;14'd11543:data <=32'h0095000B;
14'd11544:data <=32'h0091FFF2;14'd11545:data <=32'h0086FFD9;14'd11546:data <=32'h0071FFC2;
14'd11547:data <=32'h0057FFB3;14'd11548:data <=32'h0039FFAF;14'd11549:data <=32'h001CFFB5;
14'd11550:data <=32'h0004FFC4;14'd11551:data <=32'hFFF5FFDC;14'd11552:data <=32'hFFEFFFF4;
14'd11553:data <=32'hFFF2000D;14'd11554:data <=32'hFFFD0021;14'd11555:data <=32'h000E0031;
14'd11556:data <=32'h0022003C;14'd11557:data <=32'h003B0040;14'd11558:data <=32'h0056003E;
14'd11559:data <=32'h00710033;14'd11560:data <=32'h008A0020;14'd11561:data <=32'h009E0004;
14'd11562:data <=32'h00A9FFE2;14'd11563:data <=32'h00AAFFBA;14'd11564:data <=32'h009EFF96;
14'd11565:data <=32'h0088FF75;14'd11566:data <=32'h0069FF5D;14'd11567:data <=32'h0047FF51;
14'd11568:data <=32'h0026FF50;14'd11569:data <=32'h000BFF58;14'd11570:data <=32'hFFF8FF63;
14'd11571:data <=32'hFFEBFF6F;14'd11572:data <=32'hFFE4FF78;14'd11573:data <=32'hFFDFFF7D;
14'd11574:data <=32'hFFDAFF80;14'd11575:data <=32'hFFD2FF7E;14'd11576:data <=32'hFFC8FF7E;
14'd11577:data <=32'hFFBCFF7E;14'd11578:data <=32'hFFB0FF80;14'd11579:data <=32'hFFA2FF82;
14'd11580:data <=32'hFF94FF84;14'd11581:data <=32'hFF81FF88;14'd11582:data <=32'hFF6CFF8F;
14'd11583:data <=32'hFF53FF9D;14'd11584:data <=32'hFFD3FF45;14'd11585:data <=32'hFF8DFF31;
14'd11586:data <=32'hFF53FF47;14'd11587:data <=32'hFF51FFE2;14'd11588:data <=32'hFF36003B;
14'd11589:data <=32'hFF510055;14'd11590:data <=32'hFF700064;14'd11591:data <=32'hFF8D0067;
14'd11592:data <=32'hFFA30063;14'd11593:data <=32'hFFB10058;14'd11594:data <=32'hFFB60050;
14'd11595:data <=32'hFFB4004A;14'd11596:data <=32'hFFB1004B;14'd11597:data <=32'hFFAD0050;
14'd11598:data <=32'hFFAC005A;14'd11599:data <=32'hFFAD0066;14'd11600:data <=32'hFFB30074;
14'd11601:data <=32'hFFBA0083;14'd11602:data <=32'hFFC40092;14'd11603:data <=32'hFFD500A4;
14'd11604:data <=32'hFFED00B2;14'd11605:data <=32'h000C00BC;14'd11606:data <=32'h003000BE;
14'd11607:data <=32'h005700B4;14'd11608:data <=32'h007B009C;14'd11609:data <=32'h0095007A;
14'd11610:data <=32'h00A30052;14'd11611:data <=32'h00A30027;14'd11612:data <=32'h00950002;
14'd11613:data <=32'h007EFFE6;14'd11614:data <=32'h0062FFD4;14'd11615:data <=32'h0045FFCE;
14'd11616:data <=32'h002BFFCF;14'd11617:data <=32'h0015FFD8;14'd11618:data <=32'h0003FFE6;
14'd11619:data <=32'hFFF7FFF6;14'd11620:data <=32'hFFF1000A;14'd11621:data <=32'hFFF10020;
14'd11622:data <=32'hFFF70035;14'd11623:data <=32'h00050047;14'd11624:data <=32'h001B0056;
14'd11625:data <=32'h0034005E;14'd11626:data <=32'h0051005E;14'd11627:data <=32'h006B0054;
14'd11628:data <=32'h00820043;14'd11629:data <=32'h0092002E;14'd11630:data <=32'h009C0017;
14'd11631:data <=32'h00A20002;14'd11632:data <=32'h00A6FFEE;14'd11633:data <=32'h00A8FFDC;
14'd11634:data <=32'h00ABFFC8;14'd11635:data <=32'h00AFFFB1;14'd11636:data <=32'h00B0FF94;
14'd11637:data <=32'h00ACFF74;14'd11638:data <=32'h009EFF50;14'd11639:data <=32'h0088FF2D;
14'd11640:data <=32'h0065FF0F;14'd11641:data <=32'h003BFEF9;14'd11642:data <=32'h000DFEEC;
14'd11643:data <=32'hFFDEFEEB;14'd11644:data <=32'hFFB0FEF4;14'd11645:data <=32'hFF84FF04;
14'd11646:data <=32'hFF5CFF1D;14'd11647:data <=32'hFF38FF3C;14'd11648:data <=32'h003FFF7B;
14'd11649:data <=32'h001EFF44;14'd11650:data <=32'hFFDAFF23;14'd11651:data <=32'hFF1FFF78;
14'd11652:data <=32'hFEF9FFE6;14'd11653:data <=32'hFF120019;14'd11654:data <=32'hFF37003E;
14'd11655:data <=32'hFF600053;14'd11656:data <=32'hFF880056;14'd11657:data <=32'hFFA9004E;
14'd11658:data <=32'hFFBD003F;14'd11659:data <=32'hFFC8002D;14'd11660:data <=32'hFFC8001E;
14'd11661:data <=32'hFFC30013;14'd11662:data <=32'hFFBB000D;14'd11663:data <=32'hFFB0000D;
14'd11664:data <=32'hFFA50010;14'd11665:data <=32'hFF990017;14'd11666:data <=32'hFF8E0025;
14'd11667:data <=32'hFF87003A;14'd11668:data <=32'hFF850052;14'd11669:data <=32'hFF8E006E;
14'd11670:data <=32'hFFA00088;14'd11671:data <=32'hFFBB009C;14'd11672:data <=32'hFFDD00A6;
14'd11673:data <=32'hFFFE00A3;14'd11674:data <=32'h001B0098;14'd11675:data <=32'h00320085;
14'd11676:data <=32'h003F006F;14'd11677:data <=32'h0045005A;14'd11678:data <=32'h00450049;
14'd11679:data <=32'h0043003B;14'd11680:data <=32'h00400030;14'd11681:data <=32'h003D0028;
14'd11682:data <=32'h0039001F;14'd11683:data <=32'h00340017;14'd11684:data <=32'h002C0010;
14'd11685:data <=32'h0023000C;14'd11686:data <=32'h0017000A;14'd11687:data <=32'h000D000E;
14'd11688:data <=32'h00030016;14'd11689:data <=32'hFFFE0021;14'd11690:data <=32'hFFFC002E;
14'd11691:data <=32'hFFFE003A;14'd11692:data <=32'h00030048;14'd11693:data <=32'h00090054;
14'd11694:data <=32'h00140063;14'd11695:data <=32'h00220070;14'd11696:data <=32'h0036007F;
14'd11697:data <=32'h0052008C;14'd11698:data <=32'h00770092;14'd11699:data <=32'h00A2008D;
14'd11700:data <=32'h00D1007B;14'd11701:data <=32'h00FD0058;14'd11702:data <=32'h01200026;
14'd11703:data <=32'h0135FFEA;14'd11704:data <=32'h0139FFA5;14'd11705:data <=32'h012AFF63;
14'd11706:data <=32'h010CFF26;14'd11707:data <=32'h00DFFEF3;14'd11708:data <=32'h00A9FECB;
14'd11709:data <=32'h006BFEB0;14'd11710:data <=32'h002AFEA3;14'd11711:data <=32'hFFE6FEA4;
14'd11712:data <=32'h0041FF62;14'd11713:data <=32'h0030FF39;14'd11714:data <=32'h0015FF07;
14'd11715:data <=32'hFFBCFEBD;14'd11716:data <=32'hFF65FF17;14'd11717:data <=32'hFF4FFF46;
14'd11718:data <=32'hFF47FF72;14'd11719:data <=32'hFF4BFF99;14'd11720:data <=32'hFF55FFB5;
14'd11721:data <=32'hFF61FFC7;14'd11722:data <=32'hFF69FFD5;14'd11723:data <=32'hFF6FFFDF;
14'd11724:data <=32'hFF71FFE9;14'd11725:data <=32'hFF73FFF6;14'd11726:data <=32'hFF770003;
14'd11727:data <=32'hFF7D000F;14'd11728:data <=32'hFF84001A;14'd11729:data <=32'hFF8C0023;
14'd11730:data <=32'hFF940029;14'd11731:data <=32'hFF9A0030;14'd11732:data <=32'hFF9F0037;
14'd11733:data <=32'hFFA6003F;14'd11734:data <=32'hFFB00048;14'd11735:data <=32'hFFBD004E;
14'd11736:data <=32'hFFCC004F;14'd11737:data <=32'hFFDA004C;14'd11738:data <=32'hFFE50044;
14'd11739:data <=32'hFFEA0039;14'd11740:data <=32'hFFE8002E;14'd11741:data <=32'hFFE10029;
14'd11742:data <=32'hFFD8002A;14'd11743:data <=32'hFFD00031;14'd11744:data <=32'hFFCD003F;
14'd11745:data <=32'hFFD1004C;14'd11746:data <=32'hFFDC0057;14'd11747:data <=32'hFFEA005E;
14'd11748:data <=32'hFFFA005E;14'd11749:data <=32'h0008005A;14'd11750:data <=32'h00130052;
14'd11751:data <=32'h001A0047;14'd11752:data <=32'h001C003E;14'd11753:data <=32'h001A0034;
14'd11754:data <=32'h0016002C;14'd11755:data <=32'h000F0026;14'd11756:data <=32'h00050023;
14'd11757:data <=32'hFFFA0026;14'd11758:data <=32'hFFED002D;14'd11759:data <=32'hFFE1003D;
14'd11760:data <=32'hFFDA0054;14'd11761:data <=32'hFFDD0072;14'd11762:data <=32'hFFEB0093;
14'd11763:data <=32'h000700B1;14'd11764:data <=32'h003200C6;14'd11765:data <=32'h006300CE;
14'd11766:data <=32'h009800C6;14'd11767:data <=32'h00CB00AD;14'd11768:data <=32'h00F50087;
14'd11769:data <=32'h01130058;14'd11770:data <=32'h01250022;14'd11771:data <=32'h012BFFED;
14'd11772:data <=32'h0124FFB7;14'd11773:data <=32'h0116FF86;14'd11774:data <=32'h00FCFF58;
14'd11775:data <=32'h00DCFF2F;14'd11776:data <=32'h00E5FF50;14'd11777:data <=32'h00D1FF14;
14'd11778:data <=32'h00BDFEF1;14'd11779:data <=32'h00C7FF1F;14'd11780:data <=32'h007AFF42;
14'd11781:data <=32'h0064FF3C;14'd11782:data <=32'h004EFF33;14'd11783:data <=32'h003BFF2E;
14'd11784:data <=32'h0027FF23;14'd11785:data <=32'h000FFF19;14'd11786:data <=32'hFFEEFF0E;
14'd11787:data <=32'hFFC7FF0C;14'd11788:data <=32'hFF9CFF13;14'd11789:data <=32'hFF73FF28;
14'd11790:data <=32'hFF4EFF47;14'd11791:data <=32'hFF34FF6F;14'd11792:data <=32'hFF25FF9C;
14'd11793:data <=32'hFF21FFC8;14'd11794:data <=32'hFF28FFF1;14'd11795:data <=32'hFF360017;
14'd11796:data <=32'hFF4B0036;14'd11797:data <=32'hFF650050;14'd11798:data <=32'hFF840063;
14'd11799:data <=32'hFFA7006D;14'd11800:data <=32'hFFCB006E;14'd11801:data <=32'hFFEC0062;
14'd11802:data <=32'h0006004C;14'd11803:data <=32'h0016002E;14'd11804:data <=32'h00190010;
14'd11805:data <=32'h000FFFF4;14'd11806:data <=32'hFFFBFFDF;14'd11807:data <=32'hFFE2FFD7;
14'd11808:data <=32'hFFC9FFD7;14'd11809:data <=32'hFFB3FFE3;14'd11810:data <=32'hFFA5FFF3;
14'd11811:data <=32'hFF9F0006;14'd11812:data <=32'hFF9E0017;14'd11813:data <=32'hFFA00027;
14'd11814:data <=32'hFFA60034;14'd11815:data <=32'hFFAC003F;14'd11816:data <=32'hFFB40048;
14'd11817:data <=32'hFFBB004F;14'd11818:data <=32'hFFC40056;14'd11819:data <=32'hFFCD005A;
14'd11820:data <=32'hFFD6005B;14'd11821:data <=32'hFFDC005D;14'd11822:data <=32'hFFDF005D;
14'd11823:data <=32'hFFE00060;14'd11824:data <=32'hFFDF0066;14'd11825:data <=32'hFFE00070;
14'd11826:data <=32'hFFE50080;14'd11827:data <=32'hFFF20092;14'd11828:data <=32'h000500A2;
14'd11829:data <=32'h002200AB;14'd11830:data <=32'h004000AC;14'd11831:data <=32'h005F00A4;
14'd11832:data <=32'h007A0093;14'd11833:data <=32'h008D007E;14'd11834:data <=32'h00990067;
14'd11835:data <=32'h00A00051;14'd11836:data <=32'h00A50040;14'd11837:data <=32'h00A80030;
14'd11838:data <=32'h00AA0022;14'd11839:data <=32'h00B10013;14'd11840:data <=32'h01430033;
14'd11841:data <=32'h015EFFEF;14'd11842:data <=32'h014FFFB8;14'd11843:data <=32'h00C40000;
14'd11844:data <=32'h009F0027;14'd11845:data <=32'h00B3001B;14'd11846:data <=32'h00CA0007;
14'd11847:data <=32'h00DEFFEB;14'd11848:data <=32'h00EDFFC3;14'd11849:data <=32'h00F3FF92;
14'd11850:data <=32'h00E8FF5A;14'd11851:data <=32'h00CCFF25;14'd11852:data <=32'h009FFEF8;
14'd11853:data <=32'h0065FED8;14'd11854:data <=32'h0025FECD;14'd11855:data <=32'hFFE7FED1;
14'd11856:data <=32'hFFAEFEE5;14'd11857:data <=32'hFF7DFF05;14'd11858:data <=32'hFF57FF2D;
14'd11859:data <=32'hFF3DFF5A;14'd11860:data <=32'hFF2FFF8A;14'd11861:data <=32'hFF2AFFBB;
14'd11862:data <=32'hFF30FFEB;14'd11863:data <=32'hFF440016;14'd11864:data <=32'hFF630038;
14'd11865:data <=32'hFF87004F;14'd11866:data <=32'hFFAF0059;14'd11867:data <=32'hFFD60055;
14'd11868:data <=32'hFFF50045;14'd11869:data <=32'h0009002E;14'd11870:data <=32'h00130013;
14'd11871:data <=32'h0013FFFD;14'd11872:data <=32'h000CFFEA;14'd11873:data <=32'h0003FFDC;
14'd11874:data <=32'hFFF8FFD1;14'd11875:data <=32'hFFEEFFCB;14'd11876:data <=32'hFFE2FFC4;
14'd11877:data <=32'hFFD6FFBE;14'd11878:data <=32'hFFC7FFBA;14'd11879:data <=32'hFFB3FFB8;
14'd11880:data <=32'hFF9DFFBC;14'd11881:data <=32'hFF87FFC6;14'd11882:data <=32'hFF72FFD7;
14'd11883:data <=32'hFF60FFEE;14'd11884:data <=32'hFF560008;14'd11885:data <=32'hFF510025;
14'd11886:data <=32'hFF510043;14'd11887:data <=32'hFF56005F;14'd11888:data <=32'hFF5F007E;
14'd11889:data <=32'hFF6F009B;14'd11890:data <=32'hFF8600B7;14'd11891:data <=32'hFFA300D0;
14'd11892:data <=32'hFFC900E2;14'd11893:data <=32'hFFF400EA;14'd11894:data <=32'h002300E6;
14'd11895:data <=32'h004C00D5;14'd11896:data <=32'h006D00B8;14'd11897:data <=32'h00810094;
14'd11898:data <=32'h00890070;14'd11899:data <=32'h0085004F;14'd11900:data <=32'h00790038;
14'd11901:data <=32'h0067002A;14'd11902:data <=32'h00580026;14'd11903:data <=32'h004D002A;
14'd11904:data <=32'h008A00C9;14'd11905:data <=32'h00BC00BA;14'd11906:data <=32'h00DB0089;
14'd11907:data <=32'h00750026;14'd11908:data <=32'h0047005D;14'd11909:data <=32'h00590068;
14'd11910:data <=32'h0072006E;14'd11911:data <=32'h0091006C;14'd11912:data <=32'h00B3005F;
14'd11913:data <=32'h00D50043;14'd11914:data <=32'h00EE001A;14'd11915:data <=32'h00FAFFE9;
14'd11916:data <=32'h00F6FFB5;14'd11917:data <=32'h00E2FF85;14'd11918:data <=32'h00C4FF5E;
14'd11919:data <=32'h009EFF42;14'd11920:data <=32'h0077FF31;14'd11921:data <=32'h004FFF2A;
14'd11922:data <=32'h002AFF2A;14'd11923:data <=32'h0008FF30;14'd11924:data <=32'hFFE8FF3A;
14'd11925:data <=32'hFFCBFF4A;14'd11926:data <=32'hFFB2FF60;14'd11927:data <=32'hFF9FFF7A;
14'd11928:data <=32'hFF93FF97;14'd11929:data <=32'hFF92FFB3;14'd11930:data <=32'hFF97FFCC;
14'd11931:data <=32'hFFA1FFE0;14'd11932:data <=32'hFFAEFFEE;14'd11933:data <=32'hFFBAFFF7;
14'd11934:data <=32'hFFC4FFFC;14'd11935:data <=32'hFFCC0002;14'd11936:data <=32'hFFD50007;
14'd11937:data <=32'hFFE0000B;14'd11938:data <=32'hFFEF000E;14'd11939:data <=32'h0001000B;
14'd11940:data <=32'h00130002;14'd11941:data <=32'h0022FFEF;14'd11942:data <=32'h002BFFD6;
14'd11943:data <=32'h002BFFB7;14'd11944:data <=32'h001EFF99;14'd11945:data <=32'h0008FF7E;
14'd11946:data <=32'hFFE7FF6A;14'd11947:data <=32'hFFC0FF62;14'd11948:data <=32'hFF98FF62;
14'd11949:data <=32'hFF6FFF6E;14'd11950:data <=32'hFF49FF83;14'd11951:data <=32'hFF28FFA2;
14'd11952:data <=32'hFF0DFFCA;14'd11953:data <=32'hFEFAFFF8;14'd11954:data <=32'hFEF4002D;
14'd11955:data <=32'hFEFA0063;14'd11956:data <=32'hFF0E0098;14'd11957:data <=32'hFF3200C7;
14'd11958:data <=32'hFF6200E9;14'd11959:data <=32'hFF9800FC;14'd11960:data <=32'hFFCD00FD;
14'd11961:data <=32'hFFFD00F1;14'd11962:data <=32'h002100DA;14'd11963:data <=32'h003A00BD;
14'd11964:data <=32'h004600A2;14'd11965:data <=32'h004C008B;14'd11966:data <=32'h004C007B;
14'd11967:data <=32'h004A006F;14'd11968:data <=32'h00160076;14'd11969:data <=32'h001F0083;
14'd11970:data <=32'h00400088;14'd11971:data <=32'h00850079;14'd11972:data <=32'h005B009B;
14'd11973:data <=32'h006C0093;14'd11974:data <=32'h007C008A;14'd11975:data <=32'h008E007E;
14'd11976:data <=32'h00A2006E;14'd11977:data <=32'h00B40057;14'd11978:data <=32'h00C2003A;
14'd11979:data <=32'h00C80017;14'd11980:data <=32'h00C2FFF4;14'd11981:data <=32'h00B3FFD5;
14'd11982:data <=32'h009BFFBE;14'd11983:data <=32'h0082FFB0;14'd11984:data <=32'h006CFFAD;
14'd11985:data <=32'h005AFFB0;14'd11986:data <=32'h004EFFB5;14'd11987:data <=32'h0048FFB8;
14'd11988:data <=32'h0046FFBA;14'd11989:data <=32'h0043FFB8;14'd11990:data <=32'h003FFFB3;
14'd11991:data <=32'h003AFFAE;14'd11992:data <=32'h0034FFAB;14'd11993:data <=32'h002EFFA7;
14'd11994:data <=32'h0027FFA2;14'd11995:data <=32'h001FFF9E;14'd11996:data <=32'h0015FF98;
14'd11997:data <=32'h0007FF94;14'd11998:data <=32'hFFF6FF94;14'd11999:data <=32'hFFE3FF9A;
14'd12000:data <=32'hFFD2FFA6;14'd12001:data <=32'hFFC5FFBA;14'd12002:data <=32'hFFC1FFD2;
14'd12003:data <=32'hFFC7FFEB;14'd12004:data <=32'hFFD8FFFE;14'd12005:data <=32'hFFF0000A;
14'd12006:data <=32'h000A0009;14'd12007:data <=32'h0022FFFE;14'd12008:data <=32'h0035FFE8;
14'd12009:data <=32'h003EFFCD;14'd12010:data <=32'h003DFFB0;14'd12011:data <=32'h0034FF93;
14'd12012:data <=32'h0022FF7A;14'd12013:data <=32'h0009FF65;14'd12014:data <=32'hFFECFF56;
14'd12015:data <=32'hFFCAFF4E;14'd12016:data <=32'hFFA5FF4E;14'd12017:data <=32'hFF7FFF56;
14'd12018:data <=32'hFF59FF68;14'd12019:data <=32'hFF37FF84;14'd12020:data <=32'hFF1FFFAA;
14'd12021:data <=32'hFF10FFD4;14'd12022:data <=32'hFF0EFFFE;14'd12023:data <=32'hFF160025;
14'd12024:data <=32'hFF240046;14'd12025:data <=32'hFF36005E;14'd12026:data <=32'hFF470071;
14'd12027:data <=32'hFF540080;14'd12028:data <=32'hFF600091;14'd12029:data <=32'hFF6C00A2;
14'd12030:data <=32'hFF7B00B8;14'd12031:data <=32'hFF8F00CE;14'd12032:data <=32'h00150077;
14'd12033:data <=32'h00130072;14'd12034:data <=32'h0006007F;14'd12035:data <=32'hFFD50101;
14'd12036:data <=32'hFFD00134;14'd12037:data <=32'h00070137;14'd12038:data <=32'h003D0130;
14'd12039:data <=32'h0071011B;14'd12040:data <=32'h00A100FD;14'd12041:data <=32'h00CA00D7;
14'd12042:data <=32'h00E800A5;14'd12043:data <=32'h00F8006B;14'd12044:data <=32'h00F80030;
14'd12045:data <=32'h00E6FFFB;14'd12046:data <=32'h00C7FFD1;14'd12047:data <=32'h009EFFB5;
14'd12048:data <=32'h0074FFAB;14'd12049:data <=32'h004EFFAF;14'd12050:data <=32'h0033FFBD;
14'd12051:data <=32'h0022FFCF;14'd12052:data <=32'h001AFFE2;14'd12053:data <=32'h001AFFF3;
14'd12054:data <=32'h001F0000;14'd12055:data <=32'h00280009;14'd12056:data <=32'h0033000E;
14'd12057:data <=32'h003F000F;14'd12058:data <=32'h004D000B;14'd12059:data <=32'h005A0001;
14'd12060:data <=32'h0064FFF2;14'd12061:data <=32'h0067FFDF;14'd12062:data <=32'h0064FFCA;
14'd12063:data <=32'h0059FFB7;14'd12064:data <=32'h0048FFAA;14'd12065:data <=32'h0033FFA4;
14'd12066:data <=32'h0020FFA7;14'd12067:data <=32'h0011FFB0;14'd12068:data <=32'h000BFFBC;
14'd12069:data <=32'h000BFFC7;14'd12070:data <=32'h000FFFCF;14'd12071:data <=32'h0017FFD1;
14'd12072:data <=32'h001EFFCD;14'd12073:data <=32'h0022FFC6;14'd12074:data <=32'h0022FFBE;
14'd12075:data <=32'h001FFFB5;14'd12076:data <=32'h001BFFAF;14'd12077:data <=32'h0016FFAA;
14'd12078:data <=32'h0012FFA5;14'd12079:data <=32'h000EFF9F;14'd12080:data <=32'h0008FF98;
14'd12081:data <=32'h0000FF90;14'd12082:data <=32'hFFF6FF87;14'd12083:data <=32'hFFE8FF80;
14'd12084:data <=32'hFFDAFF7C;14'd12085:data <=32'hFFCAFF7A;14'd12086:data <=32'hFFBCFF7A;
14'd12087:data <=32'hFFACFF79;14'd12088:data <=32'hFF9CFF77;14'd12089:data <=32'hFF87FF75;
14'd12090:data <=32'hFF6DFF75;14'd12091:data <=32'hFF4BFF7A;14'd12092:data <=32'hFF25FF8A;
14'd12093:data <=32'hFEFEFFA8;14'd12094:data <=32'hFEDDFFD3;14'd12095:data <=32'hFEC5000C;
14'd12096:data <=32'hFF86006E;14'd12097:data <=32'hFF870077;14'd12098:data <=32'hFF79006E;
14'd12099:data <=32'hFEED0064;14'd12100:data <=32'hFECF00C6;14'd12101:data <=32'hFEFC00FD;
14'd12102:data <=32'hFF330128;14'd12103:data <=32'hFF700146;14'd12104:data <=32'hFFB40155;
14'd12105:data <=32'hFFFA0155;14'd12106:data <=32'h003E0143;14'd12107:data <=32'h00790120;
14'd12108:data <=32'h00A700EF;14'd12109:data <=32'h00C100B7;14'd12110:data <=32'h00CA007E;
14'd12111:data <=32'h00C2004C;14'd12112:data <=32'h00B00025;14'd12113:data <=32'h00970009;
14'd12114:data <=32'h007FFFF8;14'd12115:data <=32'h0069FFF0;14'd12116:data <=32'h0057FFEE;
14'd12117:data <=32'h0048FFED;14'd12118:data <=32'h003BFFEE;14'd12119:data <=32'h0031FFF1;
14'd12120:data <=32'h0026FFF6;14'd12121:data <=32'h0020FFFF;14'd12122:data <=32'h001E0008;
14'd12123:data <=32'h001F0012;14'd12124:data <=32'h00250019;14'd12125:data <=32'h002E001C;
14'd12126:data <=32'h0036001C;14'd12127:data <=32'h003C0018;14'd12128:data <=32'h00410014;
14'd12129:data <=32'h00440012;14'd12130:data <=32'h00470010;14'd12131:data <=32'h004D000F;
14'd12132:data <=32'h0055000D;14'd12133:data <=32'h00600008;14'd12134:data <=32'h006EFFFD;
14'd12135:data <=32'h0078FFEC;14'd12136:data <=32'h007CFFD6;14'd12137:data <=32'h0079FFBD;
14'd12138:data <=32'h006FFFA5;14'd12139:data <=32'h005CFF93;14'd12140:data <=32'h0045FF88;
14'd12141:data <=32'h002DFF85;14'd12142:data <=32'h0019FF89;14'd12143:data <=32'h0009FF93;
14'd12144:data <=32'h0000FF9F;14'd12145:data <=32'hFFFBFFAA;14'd12146:data <=32'hFFFBFFB3;
14'd12147:data <=32'h0000FFBA;14'd12148:data <=32'h0006FFBE;14'd12149:data <=32'h000FFFBD;
14'd12150:data <=32'h001AFFB7;14'd12151:data <=32'h0024FFAB;14'd12152:data <=32'h002BFF96;
14'd12153:data <=32'h002BFF7A;14'd12154:data <=32'h001FFF59;14'd12155:data <=32'h0006FF39;
14'd12156:data <=32'hFFDEFF1C;14'd12157:data <=32'hFFA8FF0D;14'd12158:data <=32'hFF6CFF10;
14'd12159:data <=32'hFF30FF24;14'd12160:data <=32'hFF5CFF88;14'd12161:data <=32'hFF32FF93;
14'd12162:data <=32'hFF24FF9B;14'd12163:data <=32'hFF2EFF7B;14'd12164:data <=32'hFEE3FFCC;
14'd12165:data <=32'hFEE0FFFD;14'd12166:data <=32'hFEE5002D;14'd12167:data <=32'hFEF4005A;
14'd12168:data <=32'hFF0B0083;14'd12169:data <=32'hFF2A00A8;14'd12170:data <=32'hFF5100C4;
14'd12171:data <=32'hFF7B00D4;14'd12172:data <=32'hFFA500D9;14'd12173:data <=32'hFFCA00D3;
14'd12174:data <=32'hFFE800C7;14'd12175:data <=32'hFFFD00BA;14'd12176:data <=32'h000E00AF;
14'd12177:data <=32'h001C00A5;14'd12178:data <=32'h002A009F;14'd12179:data <=32'h003C0097;
14'd12180:data <=32'h004E008D;14'd12181:data <=32'h005F007D;14'd12182:data <=32'h00700067;
14'd12183:data <=32'h0078004C;14'd12184:data <=32'h00780031;14'd12185:data <=32'h00700018;
14'd12186:data <=32'h00620003;14'd12187:data <=32'h0052FFF5;14'd12188:data <=32'h003FFFED;
14'd12189:data <=32'h002EFFEA;14'd12190:data <=32'h001BFFEC;14'd12191:data <=32'h000BFFF2;
14'd12192:data <=32'hFFFDFFFE;14'd12193:data <=32'hFFF2000E;14'd12194:data <=32'hFFED0024;
14'd12195:data <=32'hFFF1003C;14'd12196:data <=32'hFFFE0055;14'd12197:data <=32'h00150068;
14'd12198:data <=32'h00330073;14'd12199:data <=32'h00560072;14'd12200:data <=32'h00790064;
14'd12201:data <=32'h0095004C;14'd12202:data <=32'h00A7002D;14'd12203:data <=32'h00AF000A;
14'd12204:data <=32'h00ABFFE9;14'd12205:data <=32'h00A0FFCD;14'd12206:data <=32'h008FFFB8;
14'd12207:data <=32'h007DFFA9;14'd12208:data <=32'h006BFFA0;14'd12209:data <=32'h005DFF9C;
14'd12210:data <=32'h004FFF9A;14'd12211:data <=32'h0043FF99;14'd12212:data <=32'h003AFF99;
14'd12213:data <=32'h0034FF9C;14'd12214:data <=32'h0031FF9F;14'd12215:data <=32'h0032FF9F;
14'd12216:data <=32'h0037FF99;14'd12217:data <=32'h003CFF8F;14'd12218:data <=32'h003DFF7C;
14'd12219:data <=32'h0036FF64;14'd12220:data <=32'h0024FF4B;14'd12221:data <=32'h0008FF34;
14'd12222:data <=32'hFFE3FF28;14'd12223:data <=32'hFFB9FF27;14'd12224:data <=32'h0037FF1F;
14'd12225:data <=32'h0003FEF2;14'd12226:data <=32'hFFCEFEEE;14'd12227:data <=32'hFFA5FF6C;
14'd12228:data <=32'hFF64FFA5;14'd12229:data <=32'hFF65FFBA;14'd12230:data <=32'hFF6AFFCA;
14'd12231:data <=32'hFF6EFFD8;14'd12232:data <=32'hFF71FFE2;14'd12233:data <=32'hFF72FFED;
14'd12234:data <=32'hFF74FFF6;14'd12235:data <=32'hFF77FFFF;14'd12236:data <=32'hFF780004;
14'd12237:data <=32'hFF74000A;14'd12238:data <=32'hFF6E0011;14'd12239:data <=32'hFF65001D;
14'd12240:data <=32'hFF5C0030;14'd12241:data <=32'hFF56004C;14'd12242:data <=32'hFF59006E;
14'd12243:data <=32'hFF680091;14'd12244:data <=32'hFF8400B1;14'd12245:data <=32'hFFAB00C7;
14'd12246:data <=32'hFFD600D1;14'd12247:data <=32'h000300CC;14'd12248:data <=32'h002900BD;
14'd12249:data <=32'h004900A3;14'd12250:data <=32'h005F0086;14'd12251:data <=32'h006C0066;
14'd12252:data <=32'h006E0045;14'd12253:data <=32'h006B0028;14'd12254:data <=32'h0060000C;
14'd12255:data <=32'h004DFFF5;14'd12256:data <=32'h0035FFE6;14'd12257:data <=32'h0019FFDE;
14'd12258:data <=32'hFFFBFFE2;14'd12259:data <=32'hFFE1FFF1;14'd12260:data <=32'hFFCF0009;
14'd12261:data <=32'hFFC60026;14'd12262:data <=32'hFFCA0044;14'd12263:data <=32'hFFD60060;
14'd12264:data <=32'hFFED0074;14'd12265:data <=32'h00070080;14'd12266:data <=32'h00200084;
14'd12267:data <=32'h00380081;14'd12268:data <=32'h004B007B;14'd12269:data <=32'h005E0074;
14'd12270:data <=32'h006F006B;14'd12271:data <=32'h007F0063;14'd12272:data <=32'h00910059;
14'd12273:data <=32'h00A5004A;14'd12274:data <=32'h00B70037;14'd12275:data <=32'h00C6001D;
14'd12276:data <=32'h00D00000;14'd12277:data <=32'h00D5FFE1;14'd12278:data <=32'h00D4FFC1;
14'd12279:data <=32'h00CEFFA2;14'd12280:data <=32'h00C3FF83;14'd12281:data <=32'h00B5FF65;
14'd12282:data <=32'h00A2FF46;14'd12283:data <=32'h0087FF29;14'd12284:data <=32'h0063FF10;
14'd12285:data <=32'h0038FEFE;14'd12286:data <=32'h0006FEF8;14'd12287:data <=32'hFFD5FF00;
14'd12288:data <=32'h00A4FF9F;14'd12289:data <=32'h00A1FF60;14'd12290:data <=32'h0077FF27;
14'd12291:data <=32'hFFB1FF39;14'd12292:data <=32'hFF69FF80;14'd12293:data <=32'hFF6EFFA6;
14'd12294:data <=32'hFF7CFFC2;14'd12295:data <=32'hFF8FFFD6;14'd12296:data <=32'hFFA1FFE0;
14'd12297:data <=32'hFFB1FFE4;14'd12298:data <=32'hFFBFFFE2;14'd12299:data <=32'hFFCAFFDC;
14'd12300:data <=32'hFFCFFFCF;14'd12301:data <=32'hFFCDFFC1;14'd12302:data <=32'hFFC2FFB1;
14'd12303:data <=32'hFFADFFA6;14'd12304:data <=32'hFF91FFA5;14'd12305:data <=32'hFF73FFAE;
14'd12306:data <=32'hFF57FFC5;14'd12307:data <=32'hFF43FFE7;14'd12308:data <=32'hFF3B000F;
14'd12309:data <=32'hFF420038;14'd12310:data <=32'hFF54005B;14'd12311:data <=32'hFF6D0075;
14'd12312:data <=32'hFF8D0088;14'd12313:data <=32'hFFAB008F;14'd12314:data <=32'hFFC60091;
14'd12315:data <=32'hFFE0008D;14'd12316:data <=32'hFFF80086;14'd12317:data <=32'h000C007A;
14'd12318:data <=32'h001C006B;14'd12319:data <=32'h00290058;14'd12320:data <=32'h002F0043;
14'd12321:data <=32'h002F002E;14'd12322:data <=32'h0027001C;14'd12323:data <=32'h001A000E;
14'd12324:data <=32'h000A0006;14'd12325:data <=32'hFFFB0006;14'd12326:data <=32'hFFEE0009;
14'd12327:data <=32'hFFE50011;14'd12328:data <=32'hFFDD0019;14'd12329:data <=32'hFFD70021;
14'd12330:data <=32'hFFD2002A;14'd12331:data <=32'hFFCA0034;14'd12332:data <=32'hFFC40042;
14'd12333:data <=32'hFFBF0057;14'd12334:data <=32'hFFBF0071;14'd12335:data <=32'hFFC60090;
14'd12336:data <=32'hFFDA00AF;14'd12337:data <=32'hFFFA00CC;14'd12338:data <=32'h002400E0;
14'd12339:data <=32'h005600E9;14'd12340:data <=32'h008B00E4;14'd12341:data <=32'h00BE00D0;
14'd12342:data <=32'h00EC00B1;14'd12343:data <=32'h01140088;14'd12344:data <=32'h01330056;
14'd12345:data <=32'h0147001D;14'd12346:data <=32'h0150FFDF;14'd12347:data <=32'h014AFF9C;
14'd12348:data <=32'h0133FF5B;14'd12349:data <=32'h010BFF20;14'd12350:data <=32'h00D3FEF1;
14'd12351:data <=32'h0093FED3;14'd12352:data <=32'h0094FFB9;14'd12353:data <=32'h009DFF94;
14'd12354:data <=32'h00A3FF5D;14'd12355:data <=32'h0065FEEA;14'd12356:data <=32'hFFFEFF18;
14'd12357:data <=32'hFFE3FF2F;14'd12358:data <=32'hFFD0FF47;14'd12359:data <=32'hFFC6FF5D;
14'd12360:data <=32'hFFBDFF6F;14'd12361:data <=32'hFFB8FF7F;14'd12362:data <=32'hFFB5FF8F;
14'd12363:data <=32'hFFB5FF9C;14'd12364:data <=32'hFFB8FFA5;14'd12365:data <=32'hFFBBFFAB;
14'd12366:data <=32'hFFBBFFAC;14'd12367:data <=32'hFFB7FFAA;14'd12368:data <=32'hFFAEFFA8;
14'd12369:data <=32'hFFA0FFAC;14'd12370:data <=32'hFF92FFB5;14'd12371:data <=32'hFF85FFC6;
14'd12372:data <=32'hFF7FFFDB;14'd12373:data <=32'hFF7FFFF2;14'd12374:data <=32'hFF880004;
14'd12375:data <=32'hFF950011;14'd12376:data <=32'hFFA10017;14'd12377:data <=32'hFFAC0019;
14'd12378:data <=32'hFFB30018;14'd12379:data <=32'hFFB40016;14'd12380:data <=32'hFFB40018;
14'd12381:data <=32'hFFB4001D;14'd12382:data <=32'hFFB40023;14'd12383:data <=32'hFFB8002A;
14'd12384:data <=32'hFFBD0031;14'd12385:data <=32'hFFC40035;14'd12386:data <=32'hFFCA0038;
14'd12387:data <=32'hFFD1003A;14'd12388:data <=32'hFFD8003C;14'd12389:data <=32'hFFDF003D;
14'd12390:data <=32'hFFE7003B;14'd12391:data <=32'hFFF00038;14'd12392:data <=32'hFFF70030;
14'd12393:data <=32'hFFFB0024;14'd12394:data <=32'hFFFA0015;14'd12395:data <=32'hFFF00007;
14'd12396:data <=32'hFFDCFFFC;14'd12397:data <=32'hFFC3FFFB;14'd12398:data <=32'hFFA70006;
14'd12399:data <=32'hFF8E001D;14'd12400:data <=32'hFF7C003F;14'd12401:data <=32'hFF76006A;
14'd12402:data <=32'hFF7F0097;14'd12403:data <=32'hFF9600C1;14'd12404:data <=32'hFFB900E5;
14'd12405:data <=32'hFFE600FF;14'd12406:data <=32'h0017010D;14'd12407:data <=32'h004D0112;
14'd12408:data <=32'h00840109;14'd12409:data <=32'h00B800F6;14'd12410:data <=32'h00EA00D5;
14'd12411:data <=32'h011400A9;14'd12412:data <=32'h01330071;14'd12413:data <=32'h01420033;
14'd12414:data <=32'h0140FFF4;14'd12415:data <=32'h012FFFB9;14'd12416:data <=32'h0105FFDE;
14'd12417:data <=32'h0109FFAF;14'd12418:data <=32'h010EFF93;14'd12419:data <=32'h011FFFB5;
14'd12420:data <=32'h00D4FFB6;14'd12421:data <=32'h00CDFFA2;14'd12422:data <=32'h00C5FF89;
14'd12423:data <=32'h00BAFF6F;14'd12424:data <=32'h00A8FF53;14'd12425:data <=32'h008DFF3A;
14'd12426:data <=32'h006DFF26;14'd12427:data <=32'h0049FF1A;14'd12428:data <=32'h0023FF15;
14'd12429:data <=32'hFFFFFF18;14'd12430:data <=32'hFFDCFF1F;14'd12431:data <=32'hFFBBFF2D;
14'd12432:data <=32'hFF9CFF40;14'd12433:data <=32'hFF80FF5A;14'd12434:data <=32'hFF69FF79;
14'd12435:data <=32'hFF5CFFA0;14'd12436:data <=32'hFF59FFC8;14'd12437:data <=32'hFF64FFF1;
14'd12438:data <=32'hFF7B0011;14'd12439:data <=32'hFF990027;14'd12440:data <=32'hFFBB002D;
14'd12441:data <=32'hFFD80028;14'd12442:data <=32'hFFEF001A;14'd12443:data <=32'hFFFC0005;
14'd12444:data <=32'hFFFEFFF0;14'd12445:data <=32'hFFF9FFDF;14'd12446:data <=32'hFFEFFFD2;
14'd12447:data <=32'hFFE1FFCA;14'd12448:data <=32'hFFD4FFC7;14'd12449:data <=32'hFFC4FFC8;
14'd12450:data <=32'hFFB7FFCD;14'd12451:data <=32'hFFAAFFD5;14'd12452:data <=32'hFFA0FFE1;
14'd12453:data <=32'hFF99FFF0;14'd12454:data <=32'hFF970001;14'd12455:data <=32'hFF9B0011;
14'd12456:data <=32'hFFA4001D;14'd12457:data <=32'hFFAF0024;14'd12458:data <=32'hFFBA0026;
14'd12459:data <=32'hFFC30021;14'd12460:data <=32'hFFC40018;14'd12461:data <=32'hFFBE0011;
14'd12462:data <=32'hFFB1000D;14'd12463:data <=32'hFFA20012;14'd12464:data <=32'hFF920020;
14'd12465:data <=32'hFF870035;14'd12466:data <=32'hFF83004E;14'd12467:data <=32'hFF880069;
14'd12468:data <=32'hFF940081;14'd12469:data <=32'hFFA60097;14'd12470:data <=32'hFFBA00A7;
14'd12471:data <=32'hFFD000B4;14'd12472:data <=32'hFFE700BE;14'd12473:data <=32'h000000C4;
14'd12474:data <=32'h001B00C8;14'd12475:data <=32'h003800C6;14'd12476:data <=32'h005300BE;
14'd12477:data <=32'h006E00B0;14'd12478:data <=32'h0083009F;14'd12479:data <=32'h0092008B;
14'd12480:data <=32'h00FD00BF;14'd12481:data <=32'h01270093;14'd12482:data <=32'h012C006B;
14'd12483:data <=32'h00A10093;14'd12484:data <=32'h007D00AD;14'd12485:data <=32'h00A400A9;
14'd12486:data <=32'h00D00098;14'd12487:data <=32'h00FA007A;14'd12488:data <=32'h011B004C;
14'd12489:data <=32'h012F0015;14'd12490:data <=32'h0134FFD9;14'd12491:data <=32'h0128FF9D;
14'd12492:data <=32'h0111FF68;14'd12493:data <=32'h00EDFF39;14'd12494:data <=32'h00C1FF13;
14'd12495:data <=32'h008FFEF7;14'd12496:data <=32'h0056FEE7;14'd12497:data <=32'h001AFEE5;
14'd12498:data <=32'hFFDFFEF1;14'd12499:data <=32'hFFABFF0E;14'd12500:data <=32'hFF81FF37;
14'd12501:data <=32'hFF67FF69;14'd12502:data <=32'hFF5FFF9E;14'd12503:data <=32'hFF67FFCE;
14'd12504:data <=32'hFF7CFFF5;14'd12505:data <=32'hFF990010;14'd12506:data <=32'hFFB8001D;
14'd12507:data <=32'hFFD4001F;14'd12508:data <=32'hFFEC001A;14'd12509:data <=32'hFFFD0010;
14'd12510:data <=32'h000B0005;14'd12511:data <=32'h0014FFF6;14'd12512:data <=32'h001AFFE8;
14'd12513:data <=32'h001DFFD8;14'd12514:data <=32'h001AFFC7;14'd12515:data <=32'h0013FFB6;
14'd12516:data <=32'h0007FFA8;14'd12517:data <=32'hFFF7FF9C;14'd12518:data <=32'hFFE3FF96;
14'd12519:data <=32'hFFD0FF95;14'd12520:data <=32'hFFBDFF98;14'd12521:data <=32'hFFAEFF9E;
14'd12522:data <=32'hFF9FFFA4;14'd12523:data <=32'hFF90FFAC;14'd12524:data <=32'hFF81FFB4;
14'd12525:data <=32'hFF6FFFBF;14'd12526:data <=32'hFF5CFFD0;14'd12527:data <=32'hFF4CFFE8;
14'd12528:data <=32'hFF3E0005;14'd12529:data <=32'hFF3B0029;14'd12530:data <=32'hFF41004E;
14'd12531:data <=32'hFF540070;14'd12532:data <=32'hFF6E008A;14'd12533:data <=32'hFF8D009C;
14'd12534:data <=32'hFFAE00A3;14'd12535:data <=32'hFFCB00A1;14'd12536:data <=32'hFFE20099;
14'd12537:data <=32'hFFF3008E;14'd12538:data <=32'hFFFE0082;14'd12539:data <=32'h00050077;
14'd12540:data <=32'h0009006D;14'd12541:data <=32'h00080064;14'd12542:data <=32'h0004005F;
14'd12543:data <=32'hFFFD005F;14'd12544:data <=32'h000D00FA;14'd12545:data <=32'h00380104;
14'd12546:data <=32'h005900EB;14'd12547:data <=32'h000E0078;14'd12548:data <=32'hFFD700AA;
14'd12549:data <=32'hFFF200CA;14'd12550:data <=32'h001A00E1;14'd12551:data <=32'h004A00EA;
14'd12552:data <=32'h007F00E3;14'd12553:data <=32'h00AF00CD;14'd12554:data <=32'h00D700AA;
14'd12555:data <=32'h00F6007F;14'd12556:data <=32'h01080051;14'd12557:data <=32'h01100020;
14'd12558:data <=32'h010FFFF0;14'd12559:data <=32'h0104FFC1;14'd12560:data <=32'h00F0FF95;
14'd12561:data <=32'h00D0FF6D;14'd12562:data <=32'h00AAFF50;14'd12563:data <=32'h007DFF3E;
14'd12564:data <=32'h004EFF39;14'd12565:data <=32'h0024FF41;14'd12566:data <=32'h0002FF53;
14'd12567:data <=32'hFFE8FF6A;14'd12568:data <=32'hFFDBFF83;14'd12569:data <=32'hFFD4FF98;
14'd12570:data <=32'hFFD1FFAB;14'd12571:data <=32'hFFD0FFB9;14'd12572:data <=32'hFFCFFFC6;
14'd12573:data <=32'hFFCFFFD4;14'd12574:data <=32'hFFD1FFE3;14'd12575:data <=32'hFFD6FFF2;
14'd12576:data <=32'hFFE30001;14'd12577:data <=32'hFFF2000A;14'd12578:data <=32'h0008000F;
14'd12579:data <=32'h001E000A;14'd12580:data <=32'h0032FFFF;14'd12581:data <=32'h0041FFEE;
14'd12582:data <=32'h004BFFD7;14'd12583:data <=32'h004FFFBF;14'd12584:data <=32'h004CFFA2;
14'd12585:data <=32'h0043FF88;14'd12586:data <=32'h0033FF6D;14'd12587:data <=32'h001CFF54;
14'd12588:data <=32'hFFFCFF3F;14'd12589:data <=32'hFFD6FF31;14'd12590:data <=32'hFFA6FF2D;
14'd12591:data <=32'hFF75FF37;14'd12592:data <=32'hFF47FF4E;14'd12593:data <=32'hFF1FFF74;
14'd12594:data <=32'hFF03FFA7;14'd12595:data <=32'hFEF7FFDD;14'd12596:data <=32'hFEFC0013;
14'd12597:data <=32'hFF100042;14'd12598:data <=32'hFF2B0068;14'd12599:data <=32'hFF4D0081;
14'd12600:data <=32'hFF6E008F;14'd12601:data <=32'hFF8D0094;14'd12602:data <=32'hFFA90094;
14'd12603:data <=32'hFFC0008F;14'd12604:data <=32'hFFD30085;14'd12605:data <=32'hFFE00079;
14'd12606:data <=32'hFFE7006C;14'd12607:data <=32'hFFE7005F;14'd12608:data <=32'hFFB6005A;
14'd12609:data <=32'hFFAC006B;14'd12610:data <=32'hFFBB007F;14'd12611:data <=32'hFFFA0084;
14'd12612:data <=32'hFFC000A3;14'd12613:data <=32'hFFD100B6;14'd12614:data <=32'hFFED00C5;
14'd12615:data <=32'h000D00CE;14'd12616:data <=32'h003000CB;14'd12617:data <=32'h005200BE;
14'd12618:data <=32'h006C00A8;14'd12619:data <=32'h007F0090;14'd12620:data <=32'h008A0077;
14'd12621:data <=32'h00900060;14'd12622:data <=32'h0093004C;14'd12623:data <=32'h00940039;
14'd12624:data <=32'h00940028;14'd12625:data <=32'h00910015;14'd12626:data <=32'h008C0005;
14'd12627:data <=32'h0083FFF7;14'd12628:data <=32'h007AFFEC;14'd12629:data <=32'h0071FFE5;
14'd12630:data <=32'h006AFFE1;14'd12631:data <=32'h0068FFDE;14'd12632:data <=32'h0067FFD8;
14'd12633:data <=32'h0068FFCF;14'd12634:data <=32'h0065FFC0;14'd12635:data <=32'h005EFFAF;
14'd12636:data <=32'h004EFFA1;14'd12637:data <=32'h0037FF95;14'd12638:data <=32'h001FFF92;
14'd12639:data <=32'h0005FF9A;14'd12640:data <=32'hFFEFFFAB;14'd12641:data <=32'hFFE4FFC2;
14'd12642:data <=32'hFFE0FFD9;14'd12643:data <=32'hFFE6FFF1;14'd12644:data <=32'hFFF40003;
14'd12645:data <=32'h0006000F;14'd12646:data <=32'h001C0014;14'd12647:data <=32'h00340013;
14'd12648:data <=32'h004B000A;14'd12649:data <=32'h0061FFF9;14'd12650:data <=32'h0073FFE1;
14'd12651:data <=32'h007EFFC2;14'd12652:data <=32'h007FFF9D;14'd12653:data <=32'h0076FF76;
14'd12654:data <=32'h0060FF50;14'd12655:data <=32'h003FFF31;14'd12656:data <=32'h0013FF1D;
14'd12657:data <=32'hFFE4FF14;14'd12658:data <=32'hFFB5FF1C;14'd12659:data <=32'hFF8BFF2E;
14'd12660:data <=32'hFF6BFF49;14'd12661:data <=32'hFF54FF66;14'd12662:data <=32'hFF46FF83;
14'd12663:data <=32'hFF3CFF9F;14'd12664:data <=32'hFF35FFB8;14'd12665:data <=32'hFF31FFCF;
14'd12666:data <=32'hFF2CFFE7;14'd12667:data <=32'hFF2B0000;14'd12668:data <=32'hFF2C001A;
14'd12669:data <=32'hFF310034;14'd12670:data <=32'hFF3A004B;14'd12671:data <=32'hFF440061;
14'd12672:data <=32'hFFE10038;14'd12673:data <=32'hFFD10026;14'd12674:data <=32'hFFB2002B;
14'd12675:data <=32'hFF55009D;14'd12676:data <=32'hFF2E00D1;14'd12677:data <=32'hFF5700F5;
14'd12678:data <=32'hFF8A010F;14'd12679:data <=32'hFFC2011D;14'd12680:data <=32'hFFFE0119;
14'd12681:data <=32'h00350103;14'd12682:data <=32'h005F00E1;14'd12683:data <=32'h007C00B7;
14'd12684:data <=32'h0089008B;14'd12685:data <=32'h00880063;14'd12686:data <=32'h00800042;
14'd12687:data <=32'h0071002A;14'd12688:data <=32'h00600019;14'd12689:data <=32'h004E0011;
14'd12690:data <=32'h003E000C;14'd12691:data <=32'h002D000E;14'd12692:data <=32'h00200016;
14'd12693:data <=32'h00190022;14'd12694:data <=32'h00170032;14'd12695:data <=32'h00200041;
14'd12696:data <=32'h0031004D;14'd12697:data <=32'h00480050;14'd12698:data <=32'h005F004A;
14'd12699:data <=32'h00730037;14'd12700:data <=32'h0080001F;14'd12701:data <=32'h00830005;
14'd12702:data <=32'h007BFFEB;14'd12703:data <=32'h006CFFD7;14'd12704:data <=32'h005AFFCB;
14'd12705:data <=32'h0048FFC9;14'd12706:data <=32'h0037FFCA;14'd12707:data <=32'h002BFFD1;
14'd12708:data <=32'h0025FFD8;14'd12709:data <=32'h0022FFE1;14'd12710:data <=32'h0020FFE8;
14'd12711:data <=32'h0023FFEE;14'd12712:data <=32'h0028FFF5;14'd12713:data <=32'h002FFFF9;
14'd12714:data <=32'h0039FFFB;14'd12715:data <=32'h0046FFFA;14'd12716:data <=32'h0054FFF2;
14'd12717:data <=32'h005FFFE5;14'd12718:data <=32'h0067FFD3;14'd12719:data <=32'h0069FFBE;
14'd12720:data <=32'h0065FFAA;14'd12721:data <=32'h005CFF98;14'd12722:data <=32'h0051FF8A;
14'd12723:data <=32'h0046FF80;14'd12724:data <=32'h003CFF76;14'd12725:data <=32'h0035FF6B;
14'd12726:data <=32'h002DFF5D;14'd12727:data <=32'h0021FF4A;14'd12728:data <=32'h000EFF34;
14'd12729:data <=32'hFFF1FF1F;14'd12730:data <=32'hFFCCFF10;14'd12731:data <=32'hFF9DFF0B;
14'd12732:data <=32'hFF6CFF11;14'd12733:data <=32'hFF3CFF24;14'd12734:data <=32'hFF0FFF43;
14'd12735:data <=32'hFEEAFF6B;14'd12736:data <=32'hFF900012;14'd12737:data <=32'hFF8D0005;
14'd12738:data <=32'hFF76FFEA;14'd12739:data <=32'hFEDAFFB2;14'd12740:data <=32'hFE8B0003;
14'd12741:data <=32'hFE94004F;14'd12742:data <=32'hFEB20097;14'd12743:data <=32'hFEE000D4;
14'd12744:data <=32'hFF1D0101;14'd12745:data <=32'hFF630119;14'd12746:data <=32'hFFA7011C;
14'd12747:data <=32'hFFE4010E;14'd12748:data <=32'h001300F2;14'd12749:data <=32'h003500D0;
14'd12750:data <=32'h004B00AE;14'd12751:data <=32'h0057008C;14'd12752:data <=32'h005B006D;
14'd12753:data <=32'h00590052;14'd12754:data <=32'h0052003B;14'd12755:data <=32'h00450028;
14'd12756:data <=32'h0036001C;14'd12757:data <=32'h00240016;14'd12758:data <=32'h00140018;
14'd12759:data <=32'h00090021;14'd12760:data <=32'h0004002E;14'd12761:data <=32'h0006003B;
14'd12762:data <=32'h000F0044;14'd12763:data <=32'h001C0047;14'd12764:data <=32'h00270045;
14'd12765:data <=32'h002F003F;14'd12766:data <=32'h00330038;14'd12767:data <=32'h00330033;
14'd12768:data <=32'h00320031;14'd12769:data <=32'h00320033;14'd12770:data <=32'h00370036;
14'd12771:data <=32'h003F0039;14'd12772:data <=32'h004B0038;14'd12773:data <=32'h00570032;
14'd12774:data <=32'h00620028;14'd12775:data <=32'h006A001A;14'd12776:data <=32'h006C000A;
14'd12777:data <=32'h006CFFFD;14'd12778:data <=32'h0068FFF0;14'd12779:data <=32'h0062FFE7;
14'd12780:data <=32'h005BFFDE;14'd12781:data <=32'h0054FFD9;14'd12782:data <=32'h004DFFD3;
14'd12783:data <=32'h0044FFD1;14'd12784:data <=32'h003DFFD3;14'd12785:data <=32'h0036FFD7;
14'd12786:data <=32'h0033FFE0;14'd12787:data <=32'h0038FFEA;14'd12788:data <=32'h0045FFF2;
14'd12789:data <=32'h0059FFF5;14'd12790:data <=32'h0073FFEE;14'd12791:data <=32'h008FFFD8;
14'd12792:data <=32'h00A2FFB6;14'd12793:data <=32'h00ABFF89;14'd12794:data <=32'h00A4FF57;
14'd12795:data <=32'h008DFF25;14'd12796:data <=32'h0067FEFB;14'd12797:data <=32'h0036FEDB;
14'd12798:data <=32'hFFFCFEC7;14'd12799:data <=32'hFFBFFEC1;14'd12800:data <=32'hFFC2FF4F;
14'd12801:data <=32'hFFA4FF3B;14'd12802:data <=32'hFF95FF28;14'd12803:data <=32'hFF96FEEE;
14'd12804:data <=32'hFF21FF18;14'd12805:data <=32'hFEFAFF48;14'd12806:data <=32'hFEE1FF80;
14'd12807:data <=32'hFED7FFBB;14'd12808:data <=32'hFEDDFFF4;14'd12809:data <=32'hFEF10024;
14'd12810:data <=32'hFF0D0049;14'd12811:data <=32'hFF2A0063;14'd12812:data <=32'hFF480074;
14'd12813:data <=32'hFF600080;14'd12814:data <=32'hFF760088;14'd12815:data <=32'hFF8A0091;
14'd12816:data <=32'hFFA00099;14'd12817:data <=32'hFFB8009E;14'd12818:data <=32'hFFD0009E;
14'd12819:data <=32'hFFE9009A;14'd12820:data <=32'hFFFD0091;14'd12821:data <=32'h000F0083;
14'd12822:data <=32'h001C0076;14'd12823:data <=32'h00260069;14'd12824:data <=32'h002C005A;
14'd12825:data <=32'h0032004E;14'd12826:data <=32'h0036003F;14'd12827:data <=32'h0037002E;
14'd12828:data <=32'h0032001D;14'd12829:data <=32'h0028000E;14'd12830:data <=32'h00170001;
14'd12831:data <=32'h0002FFFE;14'd12832:data <=32'hFFEB0004;14'd12833:data <=32'hFFD90015;
14'd12834:data <=32'hFFCF002B;14'd12835:data <=32'hFFCF0048;14'd12836:data <=32'hFFDA0062;
14'd12837:data <=32'hFFEE0077;14'd12838:data <=32'h00080084;14'd12839:data <=32'h00240088;
14'd12840:data <=32'h003E0083;14'd12841:data <=32'h00560078;14'd12842:data <=32'h006A0067;
14'd12843:data <=32'h00790055;14'd12844:data <=32'h00830040;14'd12845:data <=32'h0088002C;
14'd12846:data <=32'h00880016;14'd12847:data <=32'h00830002;14'd12848:data <=32'h0078FFF3;
14'd12849:data <=32'h006AFFE9;14'd12850:data <=32'h005CFFE6;14'd12851:data <=32'h0051FFEB;
14'd12852:data <=32'h004BFFF5;14'd12853:data <=32'h00510000;14'd12854:data <=32'h005F0008;
14'd12855:data <=32'h00740008;14'd12856:data <=32'h008CFFFD;14'd12857:data <=32'h00A2FFE5;
14'd12858:data <=32'h00AEFFC5;14'd12859:data <=32'h00B2FFA0;14'd12860:data <=32'h00A9FF79;
14'd12861:data <=32'h0097FF57;14'd12862:data <=32'h007CFF39;14'd12863:data <=32'h005EFF22;
14'd12864:data <=32'h00B7FF52;14'd12865:data <=32'h00A6FF0E;14'd12866:data <=32'h0083FEE9;
14'd12867:data <=32'h003DFF38;14'd12868:data <=32'hFFDEFF42;14'd12869:data <=32'hFFC7FF4C;
14'd12870:data <=32'hFFB5FF5B;14'd12871:data <=32'hFFA7FF6B;14'd12872:data <=32'hFF9FFF7B;
14'd12873:data <=32'hFF9CFF88;14'd12874:data <=32'hFF9AFF8E;14'd12875:data <=32'hFF95FF8F;
14'd12876:data <=32'hFF8AFF8F;14'd12877:data <=32'hFF76FF91;14'd12878:data <=32'hFF5EFF9A;
14'd12879:data <=32'hFF46FFAE;14'd12880:data <=32'hFF32FFCB;14'd12881:data <=32'hFF25FFF0;
14'd12882:data <=32'hFF240019;14'd12883:data <=32'hFF2E0040;14'd12884:data <=32'hFF400063;
14'd12885:data <=32'hFF5A0080;14'd12886:data <=32'hFF790096;14'd12887:data <=32'hFF9B00A5;
14'd12888:data <=32'hFFBF00AB;14'd12889:data <=32'hFFE400AB;14'd12890:data <=32'h0007009F;
14'd12891:data <=32'h0027008C;14'd12892:data <=32'h0040006E;14'd12893:data <=32'h004D004A;
14'd12894:data <=32'h004D0025;14'd12895:data <=32'h003E0003;14'd12896:data <=32'h0027FFEA;
14'd12897:data <=32'h0006FFDE;14'd12898:data <=32'hFFE7FFDD;14'd12899:data <=32'hFFCCFFEA;
14'd12900:data <=32'hFFB6FFFF;14'd12901:data <=32'hFFAB0018;14'd12902:data <=32'hFFA80031;
14'd12903:data <=32'hFFAC0049;14'd12904:data <=32'hFFB6005E;14'd12905:data <=32'hFFC2006F;
14'd12906:data <=32'hFFD0007E;14'd12907:data <=32'hFFE1008B;14'd12908:data <=32'hFFF50095;
14'd12909:data <=32'h000A009C;14'd12910:data <=32'h0022009F;14'd12911:data <=32'h003B009D;
14'd12912:data <=32'h00510095;14'd12913:data <=32'h0064008B;14'd12914:data <=32'h00740080;
14'd12915:data <=32'h00830074;14'd12916:data <=32'h00910069;14'd12917:data <=32'h00A1005D;
14'd12918:data <=32'h00B3004F;14'd12919:data <=32'h00C6003B;14'd12920:data <=32'h00DA0020;
14'd12921:data <=32'h00E6FFFD;14'd12922:data <=32'h00E8FFD4;14'd12923:data <=32'h00E0FFA9;
14'd12924:data <=32'h00CBFF83;14'd12925:data <=32'h00AFFF64;14'd12926:data <=32'h008CFF51;
14'd12927:data <=32'h0068FF47;14'd12928:data <=32'h00E70019;14'd12929:data <=32'h010FFFDC;
14'd12930:data <=32'h010BFF91;14'd12931:data <=32'h0050FF58;14'd12932:data <=32'hFFF5FF6B;
14'd12933:data <=32'hFFE8FF80;14'd12934:data <=32'hFFE4FF97;14'd12935:data <=32'hFFE7FFAA;
14'd12936:data <=32'hFFF2FFB9;14'd12937:data <=32'h0003FFBF;14'd12938:data <=32'h0016FFBA;
14'd12939:data <=32'h0022FFA9;14'd12940:data <=32'h0026FF8F;14'd12941:data <=32'h001DFF73;
14'd12942:data <=32'h0005FF58;14'd12943:data <=32'hFFE3FF48;14'd12944:data <=32'hFFBCFF44;
14'd12945:data <=32'hFF93FF4D;14'd12946:data <=32'hFF6FFF63;14'd12947:data <=32'hFF53FF81;
14'd12948:data <=32'hFF3FFFA3;14'd12949:data <=32'hFF35FFC8;14'd12950:data <=32'hFF33FFED;
14'd12951:data <=32'hFF380012;14'd12952:data <=32'hFF460034;14'd12953:data <=32'hFF5B0052;
14'd12954:data <=32'hFF77006C;14'd12955:data <=32'hFF99007B;14'd12956:data <=32'hFFBD007F;
14'd12957:data <=32'hFFE00078;14'd12958:data <=32'hFFFB0067;14'd12959:data <=32'h000D0050;
14'd12960:data <=32'h00150038;14'd12961:data <=32'h00140022;14'd12962:data <=32'h000D000F;
14'd12963:data <=32'h00030003;14'd12964:data <=32'hFFF8FFFC;14'd12965:data <=32'hFFEDFFF8;
14'd12966:data <=32'hFFE4FFF6;14'd12967:data <=32'hFFD9FFF1;14'd12968:data <=32'hFFCBFFF0;
14'd12969:data <=32'hFFBBFFF1;14'd12970:data <=32'hFFA9FFF6;14'd12971:data <=32'hFF960004;
14'd12972:data <=32'hFF830019;14'd12973:data <=32'hFF770034;14'd12974:data <=32'hFF710054;
14'd12975:data <=32'hFF750077;14'd12976:data <=32'hFF7F009A;14'd12977:data <=32'hFF9400BC;
14'd12978:data <=32'hFFAF00DA;14'd12979:data <=32'hFFD100F4;14'd12980:data <=32'hFFFC0108;
14'd12981:data <=32'h002A0115;14'd12982:data <=32'h00620118;14'd12983:data <=32'h009C010E;
14'd12984:data <=32'h00D600F2;14'd12985:data <=32'h010900C8;14'd12986:data <=32'h0130008E;
14'd12987:data <=32'h0145004B;14'd12988:data <=32'h01460006;14'd12989:data <=32'h0136FFC6;
14'd12990:data <=32'h0115FF8F;14'd12991:data <=32'h00EAFF68;14'd12992:data <=32'h00960044;
14'd12993:data <=32'h00C00033;14'd12994:data <=32'h00ED0000;14'd12995:data <=32'h00DDFF6A;
14'd12996:data <=32'h0075FF62;14'd12997:data <=32'h0055FF66;14'd12998:data <=32'h003BFF70;
14'd12999:data <=32'h0028FF7E;14'd13000:data <=32'h001DFF8F;14'd13001:data <=32'h001CFF9F;
14'd13002:data <=32'h0021FFA9;14'd13003:data <=32'h002BFFAC;14'd13004:data <=32'h0032FFA3;
14'd13005:data <=32'h0034FF94;14'd13006:data <=32'h002DFF82;14'd13007:data <=32'h001EFF72;
14'd13008:data <=32'h0007FF69;14'd13009:data <=32'hFFEDFF68;14'd13010:data <=32'hFFD7FF6F;
14'd13011:data <=32'hFFC3FF7B;14'd13012:data <=32'hFFB5FF89;14'd13013:data <=32'hFFACFF97;
14'd13014:data <=32'hFFA4FFA4;14'd13015:data <=32'hFF9EFFB0;14'd13016:data <=32'hFF99FFBF;
14'd13017:data <=32'hFF95FFCD;14'd13018:data <=32'hFF95FFDC;14'd13019:data <=32'hFF97FFEA;
14'd13020:data <=32'hFF9DFFF7;14'd13021:data <=32'hFFA70001;14'd13022:data <=32'hFFAE0006;
14'd13023:data <=32'hFFB40008;14'd13024:data <=32'hFFB9000A;14'd13025:data <=32'hFFBB000D;
14'd13026:data <=32'hFFBC0011;14'd13027:data <=32'hFFC00019;14'd13028:data <=32'hFFC6001F;
14'd13029:data <=32'hFFD30025;14'd13030:data <=32'hFFE20023;14'd13031:data <=32'hFFF0001A;
14'd13032:data <=32'hFFFB000B;14'd13033:data <=32'hFFFEFFF6;14'd13034:data <=32'hFFF7FFDF;
14'd13035:data <=32'hFFE5FFCC;14'd13036:data <=32'hFFCAFFBE;14'd13037:data <=32'hFFABFFBB;
14'd13038:data <=32'hFF88FFC3;14'd13039:data <=32'hFF69FFD6;14'd13040:data <=32'hFF4EFFF1;
14'd13041:data <=32'hFF380015;14'd13042:data <=32'hFF2C003F;14'd13043:data <=32'hFF29006F;
14'd13044:data <=32'hFF3100A0;14'd13045:data <=32'hFF4700D5;14'd13046:data <=32'hFF6C0104;
14'd13047:data <=32'hFF9E012B;14'd13048:data <=32'hFFDB0144;14'd13049:data <=32'h0021014C;
14'd13050:data <=32'h00650140;14'd13051:data <=32'h00A20122;14'd13052:data <=32'h00D400F7;
14'd13053:data <=32'h00F400C4;14'd13054:data <=32'h0105008F;14'd13055:data <=32'h010C005D;
14'd13056:data <=32'h00C0006A;14'd13057:data <=32'h00DC0056;14'd13058:data <=32'h00FC004B;
14'd13059:data <=32'h011C0063;14'd13060:data <=32'h00E00040;14'd13061:data <=32'h00E30022;
14'd13062:data <=32'h00E30005;14'd13063:data <=32'h00E0FFE8;14'd13064:data <=32'h00D7FFCE;
14'd13065:data <=32'h00CCFFB6;14'd13066:data <=32'h00C1FF9F;14'd13067:data <=32'h00B4FF88;
14'd13068:data <=32'h00A3FF6E;14'd13069:data <=32'h008DFF56;14'd13070:data <=32'h006DFF41;
14'd13071:data <=32'h0047FF34;14'd13072:data <=32'h001DFF32;14'd13073:data <=32'hFFF3FF3D;
14'd13074:data <=32'hFFD1FF54;14'd13075:data <=32'hFFBAFF72;14'd13076:data <=32'hFFB0FF92;
14'd13077:data <=32'hFFAFFFB1;14'd13078:data <=32'hFFB7FFCA;14'd13079:data <=32'hFFC5FFDC;
14'd13080:data <=32'hFFD3FFE5;14'd13081:data <=32'hFFE1FFE9;14'd13082:data <=32'hFFEDFFE9;
14'd13083:data <=32'hFFF8FFE5;14'd13084:data <=32'h0000FFDE;14'd13085:data <=32'h0005FFD3;
14'd13086:data <=32'h0006FFC6;14'd13087:data <=32'h0000FFB8;14'd13088:data <=32'hFFF5FFAC;
14'd13089:data <=32'hFFE3FFA5;14'd13090:data <=32'hFFCFFFA6;14'd13091:data <=32'hFFBCFFAF;
14'd13092:data <=32'hFFAFFFBF;14'd13093:data <=32'hFFA9FFD2;14'd13094:data <=32'hFFABFFE3;
14'd13095:data <=32'hFFB4FFF1;14'd13096:data <=32'hFFC2FFF9;14'd13097:data <=32'hFFD0FFF6;
14'd13098:data <=32'hFFD8FFEE;14'd13099:data <=32'hFFDBFFE1;14'd13100:data <=32'hFFD7FFD4;
14'd13101:data <=32'hFFCBFFC9;14'd13102:data <=32'hFFBAFFC3;14'd13103:data <=32'hFFA7FFC1;
14'd13104:data <=32'hFF93FFC6;14'd13105:data <=32'hFF7EFFD0;14'd13106:data <=32'hFF6CFFDD;
14'd13107:data <=32'hFF5BFFF1;14'd13108:data <=32'hFF4C000B;14'd13109:data <=32'hFF410028;
14'd13110:data <=32'hFF3F004D;14'd13111:data <=32'hFF460071;14'd13112:data <=32'hFF560095;
14'd13113:data <=32'hFF7000B3;14'd13114:data <=32'hFF9100C8;14'd13115:data <=32'hFFB100D4;
14'd13116:data <=32'hFFD100D7;14'd13117:data <=32'hFFEB00D5;14'd13118:data <=32'h000100D2;
14'd13119:data <=32'h001400D1;14'd13120:data <=32'h0069010E;14'd13121:data <=32'h00990105;
14'd13122:data <=32'h00AD00F3;14'd13123:data <=32'h003100FC;14'd13124:data <=32'h00150102;
14'd13125:data <=32'h0043010A;14'd13126:data <=32'h00750105;14'd13127:data <=32'h00A600F4;
14'd13128:data <=32'h00D200D9;14'd13129:data <=32'h00F900B5;14'd13130:data <=32'h011B0089;
14'd13131:data <=32'h01330054;14'd13132:data <=32'h01400018;14'd13133:data <=32'h013EFFD8;
14'd13134:data <=32'h012AFF9A;14'd13135:data <=32'h0105FF60;14'd13136:data <=32'h00D2FF34;
14'd13137:data <=32'h0095FF1A;14'd13138:data <=32'h0058FF14;14'd13139:data <=32'h001FFF20;
14'd13140:data <=32'hFFF2FF3A;14'd13141:data <=32'hFFD1FF5C;14'd13142:data <=32'hFFBEFF81;
14'd13143:data <=32'hFFB6FFA3;14'd13144:data <=32'hFFB8FFC2;14'd13145:data <=32'hFFC0FFDD;
14'd13146:data <=32'hFFCEFFF2;14'd13147:data <=32'hFFDE0002;14'd13148:data <=32'hFFF3000B;
14'd13149:data <=32'h000A000F;14'd13150:data <=32'h001F000A;14'd13151:data <=32'h0032FFFC;
14'd13152:data <=32'h003DFFE9;14'd13153:data <=32'h0041FFD4;14'd13154:data <=32'h003CFFBF;
14'd13155:data <=32'h0033FFB0;14'd13156:data <=32'h0026FFA4;14'd13157:data <=32'h0019FF9E;
14'd13158:data <=32'h000DFF9C;14'd13159:data <=32'h0005FF9A;14'd13160:data <=32'hFFFEFF98;
14'd13161:data <=32'hFFF7FF90;14'd13162:data <=32'hFFEDFF89;14'd13163:data <=32'hFFDCFF81;
14'd13164:data <=32'hFFC8FF7D;14'd13165:data <=32'hFFB1FF7E;14'd13166:data <=32'hFF98FF86;
14'd13167:data <=32'hFF82FF96;14'd13168:data <=32'hFF72FFAA;14'd13169:data <=32'hFF67FFC1;
14'd13170:data <=32'hFF62FFD8;14'd13171:data <=32'hFF61FFEE;14'd13172:data <=32'hFF630002;
14'd13173:data <=32'hFF690014;14'd13174:data <=32'hFF700024;14'd13175:data <=32'hFF7A0034;
14'd13176:data <=32'hFF86003E;14'd13177:data <=32'hFF950046;14'd13178:data <=32'hFFA30047;
14'd13179:data <=32'hFFAC0043;14'd13180:data <=32'hFFAF003A;14'd13181:data <=32'hFFA90033;
14'd13182:data <=32'hFF9C0032;14'd13183:data <=32'hFF88003A;14'd13184:data <=32'hFF7900D6;
14'd13185:data <=32'hFF9300FA;14'd13186:data <=32'hFFB700F9;14'd13187:data <=32'hFF8E007F;
14'd13188:data <=32'hFF5200A0;14'd13189:data <=32'hFF6800CB;14'd13190:data <=32'hFF8A00F1;
14'd13191:data <=32'hFFB6010D;14'd13192:data <=32'hFFE7011E;14'd13193:data <=32'h001B0128;
14'd13194:data <=32'h00530123;14'd13195:data <=32'h008C0113;14'd13196:data <=32'h00C000F5;
14'd13197:data <=32'h00ED00C8;14'd13198:data <=32'h010C0092;14'd13199:data <=32'h011B0053;
14'd13200:data <=32'h01170016;14'd13201:data <=32'h0103FFE0;14'd13202:data <=32'h00E3FFB6;
14'd13203:data <=32'h00BFFF98;14'd13204:data <=32'h0098FF88;14'd13205:data <=32'h0077FF82;
14'd13206:data <=32'h0059FF82;14'd13207:data <=32'h003FFF86;14'd13208:data <=32'h0029FF8D;
14'd13209:data <=32'h0015FF95;14'd13210:data <=32'h0003FFA2;14'd13211:data <=32'hFFF5FFB2;
14'd13212:data <=32'hFFECFFC4;14'd13213:data <=32'hFFE8FFD8;14'd13214:data <=32'hFFEBFFEC;
14'd13215:data <=32'hFFF4FFFD;14'd13216:data <=32'h00010007;14'd13217:data <=32'h000F000F;
14'd13218:data <=32'h001E0011;14'd13219:data <=32'h002C0010;14'd13220:data <=32'h003A000E;
14'd13221:data <=32'h004A0008;14'd13222:data <=32'h005AFFFE;14'd13223:data <=32'h006BFFF0;
14'd13224:data <=32'h007AFFD9;14'd13225:data <=32'h0086FFBB;14'd13226:data <=32'h0086FF96;
14'd13227:data <=32'h007AFF6F;14'd13228:data <=32'h0063FF4B;14'd13229:data <=32'h003EFF2D;
14'd13230:data <=32'h0013FF1B;14'd13231:data <=32'hFFE3FF16;14'd13232:data <=32'hFFB4FF1F;
14'd13233:data <=32'hFF8CFF34;14'd13234:data <=32'hFF6AFF51;14'd13235:data <=32'hFF53FF71;
14'd13236:data <=32'hFF45FF96;14'd13237:data <=32'hFF3EFFB9;14'd13238:data <=32'hFF41FFDB;
14'd13239:data <=32'hFF48FFFB;14'd13240:data <=32'hFF590015;14'd13241:data <=32'hFF6F0027;
14'd13242:data <=32'hFF870032;14'd13243:data <=32'hFF9E0031;14'd13244:data <=32'hFFB00027;
14'd13245:data <=32'hFFB80016;14'd13246:data <=32'hFFB20005;14'd13247:data <=32'hFFA2FFF8;
14'd13248:data <=32'hFF73FFFB;14'd13249:data <=32'hFF56000D;14'd13250:data <=32'hFF55002C;
14'd13251:data <=32'hFF930040;14'd13252:data <=32'hFF4E004F;14'd13253:data <=32'hFF56006E;
14'd13254:data <=32'hFF660089;14'd13255:data <=32'hFF7D00A0;14'd13256:data <=32'hFF9400B2;
14'd13257:data <=32'hFFAE00BF;14'd13258:data <=32'hFFCA00CA;14'd13259:data <=32'hFFE900CF;
14'd13260:data <=32'h000900D0;14'd13261:data <=32'h002900C7;14'd13262:data <=32'h004600B8;
14'd13263:data <=32'h005E00A1;14'd13264:data <=32'h006D0088;14'd13265:data <=32'h00730070;
14'd13266:data <=32'h0073005C;14'd13267:data <=32'h0070004E;14'd13268:data <=32'h006E0045;
14'd13269:data <=32'h0071003E;14'd13270:data <=32'h00770036;14'd13271:data <=32'h0080002A;
14'd13272:data <=32'h00860019;14'd13273:data <=32'h00880004;14'd13274:data <=32'h0084FFED;
14'd13275:data <=32'h0077FFD9;14'd13276:data <=32'h0065FFC8;14'd13277:data <=32'h0051FFBE;
14'd13278:data <=32'h003BFFBA;14'd13279:data <=32'h0026FFBD;14'd13280:data <=32'h0015FFC5;
14'd13281:data <=32'h0005FFD1;14'd13282:data <=32'hFFFBFFE1;14'd13283:data <=32'hFFF5FFF4;
14'd13284:data <=32'hFFF50009;14'd13285:data <=32'hFFFC0020;14'd13286:data <=32'h000E0036;
14'd13287:data <=32'h00270045;14'd13288:data <=32'h004A004B;14'd13289:data <=32'h006E0044;
14'd13290:data <=32'h00920030;14'd13291:data <=32'h00AD000F;14'd13292:data <=32'h00BEFFE4;
14'd13293:data <=32'h00C0FFB6;14'd13294:data <=32'h00B5FF89;14'd13295:data <=32'h009EFF62;
14'd13296:data <=32'h007FFF44;14'd13297:data <=32'h005BFF30;14'd13298:data <=32'h0037FF25;
14'd13299:data <=32'h0013FF21;14'd13300:data <=32'hFFF2FF22;14'd13301:data <=32'hFFD2FF29;
14'd13302:data <=32'hFFB4FF35;14'd13303:data <=32'hFF99FF45;14'd13304:data <=32'hFF84FF5B;
14'd13305:data <=32'hFF74FF70;14'd13306:data <=32'hFF6BFF86;14'd13307:data <=32'hFF67FF9B;
14'd13308:data <=32'hFF66FFA9;14'd13309:data <=32'hFF64FFB5;14'd13310:data <=32'hFF5DFFBE;
14'd13311:data <=32'hFF52FFC7;14'd13312:data <=32'hFFE5FFDE;14'd13313:data <=32'hFFCDFFBF;
14'd13314:data <=32'hFFA1FFBB;14'd13315:data <=32'hFF2A0012;14'd13316:data <=32'hFEEF0034;
14'd13317:data <=32'hFF040064;14'd13318:data <=32'hFF25008B;14'd13319:data <=32'hFF4D00A9;
14'd13320:data <=32'hFF7700B7;14'd13321:data <=32'hFF9F00BA;14'd13322:data <=32'hFFC200B6;
14'd13323:data <=32'hFFE000AD;14'd13324:data <=32'hFFFA009E;14'd13325:data <=32'h000E008B;
14'd13326:data <=32'h001C0076;14'd13327:data <=32'h0022005F;14'd13328:data <=32'h001E0048;
14'd13329:data <=32'h00130038;14'd13330:data <=32'h00030030;14'd13331:data <=32'hFFF10033;
14'd13332:data <=32'hFFE60041;14'd13333:data <=32'hFFE20054;14'd13334:data <=32'hFFEA006A;
14'd13335:data <=32'hFFFB007C;14'd13336:data <=32'h00150085;14'd13337:data <=32'h00300084;
14'd13338:data <=32'h004A007A;14'd13339:data <=32'h005D0068;14'd13340:data <=32'h006B0052;
14'd13341:data <=32'h0071003C;14'd13342:data <=32'h00710026;14'd13343:data <=32'h006D0012;
14'd13344:data <=32'h00630001;14'd13345:data <=32'h0057FFF4;14'd13346:data <=32'h0048FFE9;
14'd13347:data <=32'h0036FFE5;14'd13348:data <=32'h0024FFE7;14'd13349:data <=32'h0014FFF1;
14'd13350:data <=32'h00090001;14'd13351:data <=32'h00060015;14'd13352:data <=32'h000D0028;
14'd13353:data <=32'h001C003A;14'd13354:data <=32'h00310043;14'd13355:data <=32'h00490044;
14'd13356:data <=32'h0060003D;14'd13357:data <=32'h0073002F;14'd13358:data <=32'h007F001F;
14'd13359:data <=32'h0087000D;14'd13360:data <=32'h008CFFFC;14'd13361:data <=32'h0091FFEE;
14'd13362:data <=32'h0096FFDE;14'd13363:data <=32'h009CFFCD;14'd13364:data <=32'h00A2FFB8;
14'd13365:data <=32'h00A4FF9D;14'd13366:data <=32'h00A0FF80;14'd13367:data <=32'h0095FF60;
14'd13368:data <=32'h0084FF41;14'd13369:data <=32'h006CFF25;14'd13370:data <=32'h004EFF0E;
14'd13371:data <=32'h002BFEFA;14'd13372:data <=32'h0005FEEB;14'd13373:data <=32'hFFD9FEE1;
14'd13374:data <=32'hFFA8FEDF;14'd13375:data <=32'hFF73FEE6;14'd13376:data <=32'hFFD2FFCB;
14'd13377:data <=32'hFFD0FFAF;14'd13378:data <=32'hFFBBFF86;14'd13379:data <=32'hFF28FF22;
14'd13380:data <=32'hFEBEFF4F;14'd13381:data <=32'hFEACFF99;14'd13382:data <=32'hFEAFFFE1;
14'd13383:data <=32'hFEC40025;14'd13384:data <=32'hFEE60059;14'd13385:data <=32'hFF0E0081;
14'd13386:data <=32'hFF3B009B;14'd13387:data <=32'hFF6800AA;14'd13388:data <=32'hFF9400AF;
14'd13389:data <=32'hFFBD00AA;14'd13390:data <=32'hFFE0009B;14'd13391:data <=32'hFFFC0084;
14'd13392:data <=32'h000D0067;14'd13393:data <=32'h0012004B;14'd13394:data <=32'h000C0032;
14'd13395:data <=32'hFFFC0021;14'd13396:data <=32'hFFEA001B;14'd13397:data <=32'hFFDA0020;
14'd13398:data <=32'hFFCE002C;14'd13399:data <=32'hFFCC003C;14'd13400:data <=32'hFFD1004B;
14'd13401:data <=32'hFFDB0055;14'd13402:data <=32'hFFE6005B;14'd13403:data <=32'hFFF2005D;
14'd13404:data <=32'hFFFC005B;14'd13405:data <=32'h00030059;14'd13406:data <=32'h000A0058;
14'd13407:data <=32'h00100056;14'd13408:data <=32'h00170056;14'd13409:data <=32'h001F0054;
14'd13410:data <=32'h00270050;14'd13411:data <=32'h002D004A;14'd13412:data <=32'h00320043;
14'd13413:data <=32'h0033003D;14'd13414:data <=32'h00340039;14'd13415:data <=32'h00350037;
14'd13416:data <=32'h00380036;14'd13417:data <=32'h003C0034;14'd13418:data <=32'h00410030;
14'd13419:data <=32'h0046002A;14'd13420:data <=32'h00480021;14'd13421:data <=32'h00460019;
14'd13422:data <=32'h003F0013;14'd13423:data <=32'h00360013;14'd13424:data <=32'h002E001A;
14'd13425:data <=32'h002A0028;14'd13426:data <=32'h0030003A;14'd13427:data <=32'h0041004A;
14'd13428:data <=32'h005A0056;14'd13429:data <=32'h007C0058;14'd13430:data <=32'h00A0004E;
14'd13431:data <=32'h00C30038;14'd13432:data <=32'h00E00017;14'd13433:data <=32'h00F6FFEE;
14'd13434:data <=32'h0102FFBD;14'd13435:data <=32'h0105FF88;14'd13436:data <=32'h00FBFF51;
14'd13437:data <=32'h00E3FF19;14'd13438:data <=32'h00BDFEE3;14'd13439:data <=32'h0088FEB5;
14'd13440:data <=32'h003CFF54;14'd13441:data <=32'h002DFF2D;14'd13442:data <=32'h0028FF0C;
14'd13443:data <=32'h0035FEBF;14'd13444:data <=32'hFFB2FEB9;14'd13445:data <=32'hFF7BFED9;
14'd13446:data <=32'hFF4FFF02;14'd13447:data <=32'hFF34FF31;14'd13448:data <=32'hFF24FF5E;
14'd13449:data <=32'hFF1CFF88;14'd13450:data <=32'hFF1AFFAE;14'd13451:data <=32'hFF1EFFD1;
14'd13452:data <=32'hFF26FFF2;14'd13453:data <=32'hFF340011;14'd13454:data <=32'hFF46002A;
14'd13455:data <=32'hFF5B003D;14'd13456:data <=32'hFF73004A;14'd13457:data <=32'hFF87004F;
14'd13458:data <=32'hFF980050;14'd13459:data <=32'hFFA50051;14'd13460:data <=32'hFFAF0052;
14'd13461:data <=32'hFFB70056;14'd13462:data <=32'hFFC2005B;14'd13463:data <=32'hFFD1005E;
14'd13464:data <=32'hFFE3005D;14'd13465:data <=32'hFFF50057;14'd13466:data <=32'h00030049;
14'd13467:data <=32'h000B0036;14'd13468:data <=32'h000A0023;14'd13469:data <=32'h00010013;
14'd13470:data <=32'hFFF20009;14'd13471:data <=32'hFFE10007;14'd13472:data <=32'hFFD0000C;
14'd13473:data <=32'hFFC40019;14'd13474:data <=32'hFFBC0028;14'd13475:data <=32'hFFBA0038;
14'd13476:data <=32'hFFBD004A;14'd13477:data <=32'hFFC3005B;14'd13478:data <=32'hFFCE006B;
14'd13479:data <=32'hFFDD0078;14'd13480:data <=32'hFFF00082;14'd13481:data <=32'h00070086;
14'd13482:data <=32'h001E0084;14'd13483:data <=32'h0035007C;14'd13484:data <=32'h0047006C;
14'd13485:data <=32'h00530056;14'd13486:data <=32'h00530041;14'd13487:data <=32'h004C002E;
14'd13488:data <=32'h003E0024;14'd13489:data <=32'h002E0023;14'd13490:data <=32'h0022002D;
14'd13491:data <=32'h001D003E;14'd13492:data <=32'h00220052;14'd13493:data <=32'h00310064;
14'd13494:data <=32'h00480071;14'd13495:data <=32'h00660075;14'd13496:data <=32'h00850071;
14'd13497:data <=32'h00A50063;14'd13498:data <=32'h00C2004F;14'd13499:data <=32'h00DA0033;
14'd13500:data <=32'h00F0000F;14'd13501:data <=32'h00FEFFE5;14'd13502:data <=32'h0103FFB6;
14'd13503:data <=32'h00FCFF83;14'd13504:data <=32'h0112FFC3;14'd13505:data <=32'h0121FF79;
14'd13506:data <=32'h0114FF47;14'd13507:data <=32'h00C7FF71;14'd13508:data <=32'h0069FF4D;
14'd13509:data <=32'h004FFF4B;14'd13510:data <=32'h003AFF4E;14'd13511:data <=32'h002BFF50;
14'd13512:data <=32'h0020FF50;14'd13513:data <=32'h0015FF4A;14'd13514:data <=32'h0004FF42;
14'd13515:data <=32'hFFF0FF3A;14'd13516:data <=32'hFFD4FF36;14'd13517:data <=32'hFFB6FF39;
14'd13518:data <=32'hFF98FF43;14'd13519:data <=32'hFF7CFF54;14'd13520:data <=32'hFF63FF69;
14'd13521:data <=32'hFF4FFF83;14'd13522:data <=32'hFF3EFF9F;14'd13523:data <=32'hFF31FFC0;
14'd13524:data <=32'hFF2BFFE5;14'd13525:data <=32'hFF2D000D;14'd13526:data <=32'hFF390035;
14'd13527:data <=32'hFF51005B;14'd13528:data <=32'hFF730077;14'd13529:data <=32'hFF9F0087;
14'd13530:data <=32'hFFC90087;14'd13531:data <=32'hFFF2007A;14'd13532:data <=32'h000E0062;
14'd13533:data <=32'h00210042;14'd13534:data <=32'h00250022;14'd13535:data <=32'h001E0004;
14'd13536:data <=32'h0010FFEE;14'd13537:data <=32'hFFFCFFDF;14'd13538:data <=32'hFFE6FFD7;
14'd13539:data <=32'hFFCFFFD7;14'd13540:data <=32'hFFB9FFDD;14'd13541:data <=32'hFFA5FFE8;
14'd13542:data <=32'hFF96FFF8;14'd13543:data <=32'hFF89000E;14'd13544:data <=32'hFF830027;
14'd13545:data <=32'hFF840042;14'd13546:data <=32'hFF8D005C;14'd13547:data <=32'hFF9D0071;
14'd13548:data <=32'hFFB10081;14'd13549:data <=32'hFFC50089;14'd13550:data <=32'hFFD8008B;
14'd13551:data <=32'hFFE7008B;14'd13552:data <=32'hFFF1008A;14'd13553:data <=32'hFFF9008D;
14'd13554:data <=32'h00010093;14'd13555:data <=32'h000E009C;14'd13556:data <=32'h002000A5;
14'd13557:data <=32'h003800AB;14'd13558:data <=32'h005600AB;14'd13559:data <=32'h007300A2;
14'd13560:data <=32'h008E0091;14'd13561:data <=32'h00A5007A;14'd13562:data <=32'h00B50061;
14'd13563:data <=32'h00C00045;14'd13564:data <=32'h00C5002A;14'd13565:data <=32'h00C8000F;
14'd13566:data <=32'h00C6FFF4;14'd13567:data <=32'h00C0FFDA;14'd13568:data <=32'h00E200AC;
14'd13569:data <=32'h0127007F;14'd13570:data <=32'h01400035;14'd13571:data <=32'h00A3FFC4;
14'd13572:data <=32'h004DFFB0;14'd13573:data <=32'h0040FFC0;14'd13574:data <=32'h003FFFD2;
14'd13575:data <=32'h0047FFE1;14'd13576:data <=32'h005AFFE7;14'd13577:data <=32'h0070FFE1;
14'd13578:data <=32'h0083FFCD;14'd13579:data <=32'h008FFFB0;14'd13580:data <=32'h008EFF8E;
14'd13581:data <=32'h0082FF6D;14'd13582:data <=32'h006DFF4E;14'd13583:data <=32'h0050FF35;
14'd13584:data <=32'h002DFF23;14'd13585:data <=32'h0006FF1A;14'd13586:data <=32'hFFDCFF17;
14'd13587:data <=32'hFFB1FF1F;14'd13588:data <=32'hFF86FF31;14'd13589:data <=32'hFF60FF4F;
14'd13590:data <=32'hFF43FF78;14'd13591:data <=32'hFF34FFA7;14'd13592:data <=32'hFF33FFD9;
14'd13593:data <=32'hFF410007;14'd13594:data <=32'hFF5B002B;14'd13595:data <=32'hFF7D0042;
14'd13596:data <=32'hFFA0004E;14'd13597:data <=32'hFFBF004D;14'd13598:data <=32'hFFD90045;
14'd13599:data <=32'hFFEC0038;14'd13600:data <=32'hFFF90029;14'd13601:data <=32'h0002001A;
14'd13602:data <=32'h0007000B;14'd13603:data <=32'h0009FFFA;14'd13604:data <=32'h0007FFEA;
14'd13605:data <=32'h0000FFD9;14'd13606:data <=32'hFFF4FFCA;14'd13607:data <=32'hFFE2FFBD;
14'd13608:data <=32'hFFCCFFB7;14'd13609:data <=32'hFFB5FFB9;14'd13610:data <=32'hFF9DFFBE;
14'd13611:data <=32'hFF89FFCA;14'd13612:data <=32'hFF75FFDA;14'd13613:data <=32'hFF64FFED;
14'd13614:data <=32'hFF560002;14'd13615:data <=32'hFF4A001C;14'd13616:data <=32'hFF40003A;
14'd13617:data <=32'hFF39005F;14'd13618:data <=32'hFF3C0089;14'd13619:data <=32'hFF4B00B7;
14'd13620:data <=32'hFF6600E5;14'd13621:data <=32'hFF90010A;14'd13622:data <=32'hFFC60125;
14'd13623:data <=32'h00020131;14'd13624:data <=32'h003F012A;14'd13625:data <=32'h00770115;
14'd13626:data <=32'h00A600F4;14'd13627:data <=32'h00CA00CB;14'd13628:data <=32'h00E2009C;
14'd13629:data <=32'h00EF006D;14'd13630:data <=32'h00F2003F;14'd13631:data <=32'h00E90013;
14'd13632:data <=32'h004E00B9;14'd13633:data <=32'h008400BD;14'd13634:data <=32'h00C5009E;
14'd13635:data <=32'h00E5FFFC;14'd13636:data <=32'h0088FFD0;14'd13637:data <=32'h006DFFD2;
14'd13638:data <=32'h005AFFDC;14'd13639:data <=32'h0051FFEC;14'd13640:data <=32'h0054FFFA;
14'd13641:data <=32'h00600003;14'd13642:data <=32'h00710000;14'd13643:data <=32'h0080FFF4;
14'd13644:data <=32'h008AFFE2;14'd13645:data <=32'h008EFFCB;14'd13646:data <=32'h008CFFB4;
14'd13647:data <=32'h0082FF9F;14'd13648:data <=32'h0076FF8B;14'd13649:data <=32'h0067FF7B;
14'd13650:data <=32'h0054FF6B;14'd13651:data <=32'h003DFF5E;14'd13652:data <=32'h0023FF55;
14'd13653:data <=32'h0006FF55;14'd13654:data <=32'hFFE8FF5A;14'd13655:data <=32'hFFCFFF69;
14'd13656:data <=32'hFFBBFF7D;14'd13657:data <=32'hFFB0FF94;14'd13658:data <=32'hFFADFFAA;
14'd13659:data <=32'hFFAFFFBC;14'd13660:data <=32'hFFB3FFC8;14'd13661:data <=32'hFFB7FFCF;
14'd13662:data <=32'hFFB9FFD7;14'd13663:data <=32'hFFB8FFDC;14'd13664:data <=32'hFFB8FFE5;
14'd13665:data <=32'hFFB9FFF0;14'd13666:data <=32'hFFBEFFFC;14'd13667:data <=32'hFFCA0007;
14'd13668:data <=32'hFFD9000F;14'd13669:data <=32'hFFEA000E;14'd13670:data <=32'hFFFC0007;
14'd13671:data <=32'h0009FFF8;14'd13672:data <=32'h0010FFE5;14'd13673:data <=32'h0013FFCF;
14'd13674:data <=32'h000DFFBA;14'd13675:data <=32'h0000FFA4;14'd13676:data <=32'hFFEDFF92;
14'd13677:data <=32'hFFD4FF81;14'd13678:data <=32'hFFB4FF76;14'd13679:data <=32'hFF8EFF73;
14'd13680:data <=32'hFF63FF7B;14'd13681:data <=32'hFF35FF8E;14'd13682:data <=32'hFF0CFFB3;
14'd13683:data <=32'hFEEBFFE4;14'd13684:data <=32'hFED90021;14'd13685:data <=32'hFED90065;
14'd13686:data <=32'hFEEC00A6;14'd13687:data <=32'hFF1100DE;14'd13688:data <=32'hFF43010C;
14'd13689:data <=32'hFF7C0128;14'd13690:data <=32'hFFB80135;14'd13691:data <=32'hFFF10134;
14'd13692:data <=32'h00250129;14'd13693:data <=32'h00540113;14'd13694:data <=32'h007C00F9;
14'd13695:data <=32'h009C00D7;14'd13696:data <=32'h004A00B7;14'd13697:data <=32'h006A00B7;
14'd13698:data <=32'h008E00BD;14'd13699:data <=32'h00B800D6;14'd13700:data <=32'h0087009E;
14'd13701:data <=32'h0090008C;14'd13702:data <=32'h0099007E;14'd13703:data <=32'h00A10070;
14'd13704:data <=32'h00B10062;14'd13705:data <=32'h00BF004E;14'd13706:data <=32'h00CE0034;
14'd13707:data <=32'h00D60013;14'd13708:data <=32'h00D3FFED;14'd13709:data <=32'h00C8FFCB;
14'd13710:data <=32'h00B2FFAC;14'd13711:data <=32'h0098FF95;14'd13712:data <=32'h007AFF89;
14'd13713:data <=32'h005FFF85;14'd13714:data <=32'h0047FF85;14'd13715:data <=32'h0031FF8B;
14'd13716:data <=32'h0020FF93;14'd13717:data <=32'h0011FF9D;14'd13718:data <=32'h0006FFAA;
14'd13719:data <=32'hFFFEFFBA;14'd13720:data <=32'hFFFEFFC8;14'd13721:data <=32'h0003FFD5;
14'd13722:data <=32'h000EFFDE;14'd13723:data <=32'h001CFFDE;14'd13724:data <=32'h0028FFD6;
14'd13725:data <=32'h002FFFC8;14'd13726:data <=32'h002DFFB7;14'd13727:data <=32'h0024FFA6;
14'd13728:data <=32'h0013FF9B;14'd13729:data <=32'hFFFFFF9A;14'd13730:data <=32'hFFEBFF9F;
14'd13731:data <=32'hFFDDFFA9;14'd13732:data <=32'hFFD5FFBA;14'd13733:data <=32'hFFD4FFC9;
14'd13734:data <=32'hFFD9FFD5;14'd13735:data <=32'hFFE2FFE0;14'd13736:data <=32'hFFECFFE1;
14'd13737:data <=32'hFFF7FFE0;14'd13738:data <=32'h0001FFD9;14'd13739:data <=32'h0008FFCE;
14'd13740:data <=32'h000CFFC0;14'd13741:data <=32'h000CFFB0;14'd13742:data <=32'h0006FF9A;
14'd13743:data <=32'hFFF7FF85;14'd13744:data <=32'hFFE1FF73;14'd13745:data <=32'hFFC1FF65;
14'd13746:data <=32'hFF9AFF63;14'd13747:data <=32'hFF72FF6B;14'd13748:data <=32'hFF4CFF81;
14'd13749:data <=32'hFF2EFFA2;14'd13750:data <=32'hFF1AFFCB;14'd13751:data <=32'hFF11FFF4;
14'd13752:data <=32'hFF14001D;14'd13753:data <=32'hFF1E003E;14'd13754:data <=32'hFF2C005C;
14'd13755:data <=32'hFF3A0075;14'd13756:data <=32'hFF49008C;14'd13757:data <=32'hFF5A00A2;
14'd13758:data <=32'hFF6E00B7;14'd13759:data <=32'hFF8500CB;14'd13760:data <=32'hFFD4010B;
14'd13761:data <=32'hFFFF0114;14'd13762:data <=32'h0015010D;14'd13763:data <=32'hFFA100F9;
14'd13764:data <=32'hFF8100F1;14'd13765:data <=32'hFFA4010D;14'd13766:data <=32'hFFCE0125;
14'd13767:data <=32'hFFFD0133;14'd13768:data <=32'h00360139;14'd13769:data <=32'h00740130;
14'd13770:data <=32'h00B10117;14'd13771:data <=32'h00E500EC;14'd13772:data <=32'h010D00B3;
14'd13773:data <=32'h01210072;14'd13774:data <=32'h0123002F;14'd13775:data <=32'h0113FFF4;
14'd13776:data <=32'h00F6FFC1;14'd13777:data <=32'h00D1FF9C;14'd13778:data <=32'h00A8FF84;
14'd13779:data <=32'h007EFF78;14'd13780:data <=32'h0056FF75;14'd13781:data <=32'h0031FF7C;
14'd13782:data <=32'h0010FF8B;14'd13783:data <=32'hFFF7FFA2;14'd13784:data <=32'hFFE7FFBE;
14'd13785:data <=32'hFFE2FFDD;14'd13786:data <=32'hFFE9FFF9;14'd13787:data <=32'hFFFA000E;
14'd13788:data <=32'h0011001B;14'd13789:data <=32'h0029001C;14'd13790:data <=32'h003F0013;
14'd13791:data <=32'h004D0004;14'd13792:data <=32'h0054FFF2;14'd13793:data <=32'h0054FFE1;
14'd13794:data <=32'h004FFFD4;14'd13795:data <=32'h0048FFCB;14'd13796:data <=32'h0043FFC5;
14'd13797:data <=32'h003FFFC0;14'd13798:data <=32'h003DFFBA;14'd13799:data <=32'h003BFFB3;
14'd13800:data <=32'h0037FFAA;14'd13801:data <=32'h0031FF9F;14'd13802:data <=32'h0029FF96;
14'd13803:data <=32'h001DFF90;14'd13804:data <=32'h0011FF89;14'd13805:data <=32'h0006FF86;
14'd13806:data <=32'hFFFBFF83;14'd13807:data <=32'hFFEFFF80;14'd13808:data <=32'hFFE1FF7F;
14'd13809:data <=32'hFFD1FF7E;14'd13810:data <=32'hFFBEFF80;14'd13811:data <=32'hFFADFF88;
14'd13812:data <=32'hFF9CFF95;14'd13813:data <=32'hFF90FFA5;14'd13814:data <=32'hFF8BFFB7;
14'd13815:data <=32'hFF8DFFC8;14'd13816:data <=32'hFF93FFD1;14'd13817:data <=32'hFF9AFFD4;
14'd13818:data <=32'hFF9CFFD2;14'd13819:data <=32'hFF97FFCA;14'd13820:data <=32'hFF8AFFC2;
14'd13821:data <=32'hFF75FFC2;14'd13822:data <=32'hFF5BFFC8;14'd13823:data <=32'hFF3FFFDB;
14'd13824:data <=32'hFF1A0078;14'd13825:data <=32'hFF26009F;14'd13826:data <=32'hFF4400A5;
14'd13827:data <=32'hFF39001F;14'd13828:data <=32'hFEF00025;14'd13829:data <=32'hFEEA005B;
14'd13830:data <=32'hFEF20094;14'd13831:data <=32'hFF0700CE;14'd13832:data <=32'hFF2D0104;
14'd13833:data <=32'hFF630130;14'd13834:data <=32'hFFA6014C;14'd13835:data <=32'hFFF00154;
14'd13836:data <=32'h00370147;14'd13837:data <=32'h00730129;14'd13838:data <=32'h00A400FE;
14'd13839:data <=32'h00C300CC;14'd13840:data <=32'h00D50099;14'd13841:data <=32'h00DB0068;
14'd13842:data <=32'h00D6003C;14'd13843:data <=32'h00CA0017;14'd13844:data <=32'h00BAFFF5;
14'd13845:data <=32'h00A3FFD9;14'd13846:data <=32'h0088FFC3;14'd13847:data <=32'h006AFFB7;
14'd13848:data <=32'h004BFFB4;14'd13849:data <=32'h0030FFB9;14'd13850:data <=32'h001AFFC6;
14'd13851:data <=32'h000CFFD7;14'd13852:data <=32'h0007FFE7;14'd13853:data <=32'h0006FFF6;
14'd13854:data <=32'h000A0002;14'd13855:data <=32'h000D0008;14'd13856:data <=32'h00100010;
14'd13857:data <=32'h00140018;14'd13858:data <=32'h00180020;14'd13859:data <=32'h0022002B;
14'd13860:data <=32'h00310034;14'd13861:data <=32'h00460039;14'd13862:data <=32'h005E0038;
14'd13863:data <=32'h0079002C;14'd13864:data <=32'h00900018;14'd13865:data <=32'h00A1FFFB;
14'd13866:data <=32'h00A9FFD8;14'd13867:data <=32'h00A8FFB6;14'd13868:data <=32'h009DFF92;
14'd13869:data <=32'h008BFF75;14'd13870:data <=32'h0073FF5B;14'd13871:data <=32'h0056FF48;
14'd13872:data <=32'h0035FF3C;14'd13873:data <=32'h0012FF36;14'd13874:data <=32'hFFF0FF38;
14'd13875:data <=32'hFFCDFF43;14'd13876:data <=32'hFFB0FF57;14'd13877:data <=32'hFF9AFF73;
14'd13878:data <=32'hFF8FFF93;14'd13879:data <=32'hFF91FFB2;14'd13880:data <=32'hFF9EFFC9;
14'd13881:data <=32'hFFB1FFD8;14'd13882:data <=32'hFFC6FFD8;14'd13883:data <=32'hFFD6FFCD;
14'd13884:data <=32'hFFDCFFB9;14'd13885:data <=32'hFFD6FFA5;14'd13886:data <=32'hFFC5FF92;
14'd13887:data <=32'hFFABFF86;14'd13888:data <=32'hFF78FF98;14'd13889:data <=32'hFF58FF9D;
14'd13890:data <=32'hFF51FFB4;14'd13891:data <=32'hFF8CFFC7;14'd13892:data <=32'hFF3DFFB1;
14'd13893:data <=32'hFF29FFCD;14'd13894:data <=32'hFF18FFEF;14'd13895:data <=32'hFF110016;
14'd13896:data <=32'hFF120041;14'd13897:data <=32'hFF1F006E;14'd13898:data <=32'hFF390094;
14'd13899:data <=32'hFF5C00B1;14'd13900:data <=32'hFF8400C2;14'd13901:data <=32'hFFA900C8;
14'd13902:data <=32'hFFCB00C4;14'd13903:data <=32'hFFE600BB;14'd13904:data <=32'hFFFA00B1;
14'd13905:data <=32'h000B00A9;14'd13906:data <=32'h001900A3;14'd13907:data <=32'h002A009C;
14'd13908:data <=32'h003A0094;14'd13909:data <=32'h004C0088;14'd13910:data <=32'h005B0077;
14'd13911:data <=32'h00650064;14'd13912:data <=32'h006D0050;14'd13913:data <=32'h006E003C;
14'd13914:data <=32'h006C002A;14'd13915:data <=32'h0068001A;14'd13916:data <=32'h00630009;
14'd13917:data <=32'h005AFFFB;14'd13918:data <=32'h004FFFEC;14'd13919:data <=32'h003EFFE1;
14'd13920:data <=32'h0029FFDA;14'd13921:data <=32'h0011FFDB;14'd13922:data <=32'hFFF9FFE7;
14'd13923:data <=32'hFFE6FFFD;14'd13924:data <=32'hFFDD0019;14'd13925:data <=32'hFFDF003B;
14'd13926:data <=32'hFFEF0059;14'd13927:data <=32'h000B0071;14'd13928:data <=32'h002E007F;
14'd13929:data <=32'h00560080;14'd13930:data <=32'h007B0074;14'd13931:data <=32'h009B005F;
14'd13932:data <=32'h00B50042;14'd13933:data <=32'h00C70020;14'd13934:data <=32'h00D1FFFB;
14'd13935:data <=32'h00D2FFD4;14'd13936:data <=32'h00CCFFAE;14'd13937:data <=32'h00BDFF8B;
14'd13938:data <=32'h00A6FF6A;14'd13939:data <=32'h0087FF50;14'd13940:data <=32'h0065FF41;
14'd13941:data <=32'h0041FF3C;14'd13942:data <=32'h0020FF41;14'd13943:data <=32'h0006FF4C;
14'd13944:data <=32'hFFF7FF5B;14'd13945:data <=32'hFFEEFF67;14'd13946:data <=32'hFFEBFF6E;
14'd13947:data <=32'hFFE7FF6E;14'd13948:data <=32'hFFE1FF69;14'd13949:data <=32'hFFD4FF62;
14'd13950:data <=32'hFFC1FF5E;14'd13951:data <=32'hFFA9FF5E;14'd13952:data <=32'h001BFFAF;
14'd13953:data <=32'h0014FF87;14'd13954:data <=32'hFFF3FF71;14'd13955:data <=32'hFF73FF9B;
14'd13956:data <=32'hFF2EFF92;14'd13957:data <=32'hFF27FFB6;14'd13958:data <=32'hFF26FFD9;
14'd13959:data <=32'hFF2CFFFB;14'd13960:data <=32'hFF38001C;14'd13961:data <=32'hFF4A0039;
14'd13962:data <=32'hFF64004F;14'd13963:data <=32'hFF82005C;14'd13964:data <=32'hFF9F005D;
14'd13965:data <=32'hFFB80056;14'd13966:data <=32'hFFC70047;14'd13967:data <=32'hFFCD0035;
14'd13968:data <=32'hFFC60028;14'd13969:data <=32'hFFB90023;14'd13970:data <=32'hFFAC0027;
14'd13971:data <=32'hFFA10035;14'd13972:data <=32'hFF9D0049;14'd13973:data <=32'hFFA2005F;
14'd13974:data <=32'hFFAD0073;14'd13975:data <=32'hFFBD0081;14'd13976:data <=32'hFFD2008D;
14'd13977:data <=32'hFFE80092;14'd13978:data <=32'h00010094;14'd13979:data <=32'h00190091;
14'd13980:data <=32'h00310086;14'd13981:data <=32'h00480076;14'd13982:data <=32'h0059005E;
14'd13983:data <=32'h00610042;14'd13984:data <=32'h00600026;14'd13985:data <=32'h0053000B;
14'd13986:data <=32'h003FFFF7;14'd13987:data <=32'h0025FFEE;14'd13988:data <=32'h0009FFF1;
14'd13989:data <=32'hFFF3FFFF;14'd13990:data <=32'hFFE50013;14'd13991:data <=32'hFFE1002B;
14'd13992:data <=32'hFFE60042;14'd13993:data <=32'hFFF10056;14'd13994:data <=32'h00020064;
14'd13995:data <=32'h0014006E;14'd13996:data <=32'h00280073;14'd13997:data <=32'h003C0075;
14'd13998:data <=32'h00500075;14'd13999:data <=32'h00670071;14'd14000:data <=32'h007D006A;
14'd14001:data <=32'h0094005C;14'd14002:data <=32'h00A80049;14'd14003:data <=32'h00BA0033;
14'd14004:data <=32'h00C60019;14'd14005:data <=32'h00CDFFFE;14'd14006:data <=32'h00D0FFE4;
14'd14007:data <=32'h00D2FFC9;14'd14008:data <=32'h00D3FFAE;14'd14009:data <=32'h00D2FF8F;
14'd14010:data <=32'h00CCFF6D;14'd14011:data <=32'h00C0FF46;14'd14012:data <=32'h00A9FF1D;
14'd14013:data <=32'h0084FEF5;14'd14014:data <=32'h0054FED8;14'd14015:data <=32'h001BFEC6;
14'd14016:data <=32'h001CFFCD;14'd14017:data <=32'h0030FFB3;14'd14018:data <=32'h0034FF81;
14'd14019:data <=32'hFFC8FEEB;14'd14020:data <=32'hFF5FFEE2;14'd14021:data <=32'hFF35FF10;
14'd14022:data <=32'hFF18FF43;14'd14023:data <=32'hFF09FF7A;14'd14024:data <=32'hFF06FFB1;
14'd14025:data <=32'hFF0EFFE5;14'd14026:data <=32'hFF260013;14'd14027:data <=32'hFF480037;
14'd14028:data <=32'hFF70004B;14'd14029:data <=32'hFF990050;14'd14030:data <=32'hFFBB0047;
14'd14031:data <=32'hFFD20034;14'd14032:data <=32'hFFDD001C;14'd14033:data <=32'hFFDB0007;
14'd14034:data <=32'hFFCFFFF8;14'd14035:data <=32'hFFC0FFF4;14'd14036:data <=32'hFFB1FFF6;
14'd14037:data <=32'hFFA6FFFF;14'd14038:data <=32'hFF9F000C;14'd14039:data <=32'hFF9A0019;
14'd14040:data <=32'hFF9A0028;14'd14041:data <=32'hFF9D0036;14'd14042:data <=32'hFFA10043;
14'd14043:data <=32'hFFAB0052;14'd14044:data <=32'hFFB7005E;14'd14045:data <=32'hFFC70068;
14'd14046:data <=32'hFFDA006C;14'd14047:data <=32'hFFED006A;14'd14048:data <=32'hFFFD0062;
14'd14049:data <=32'h00080056;14'd14050:data <=32'h000C004A;14'd14051:data <=32'h000B0040;
14'd14052:data <=32'h0007003A;14'd14053:data <=32'h00030039;14'd14054:data <=32'h0001003C;
14'd14055:data <=32'h0002003F;14'd14056:data <=32'h00060040;14'd14057:data <=32'h000D003F;
14'd14058:data <=32'h000F003B;14'd14059:data <=32'h000E0034;14'd14060:data <=32'h000A0030;
14'd14061:data <=32'h00020030;14'd14062:data <=32'hFFF80035;14'd14063:data <=32'hFFF00042;
14'd14064:data <=32'hFFED0054;14'd14065:data <=32'hFFF10068;14'd14066:data <=32'hFFFD007E;
14'd14067:data <=32'h00100091;14'd14068:data <=32'h002900A1;14'd14069:data <=32'h004800AC;
14'd14070:data <=32'h006B00B2;14'd14071:data <=32'h009400B0;14'd14072:data <=32'h00C100A6;
14'd14073:data <=32'h00EF008F;14'd14074:data <=32'h011C0068;14'd14075:data <=32'h01410033;
14'd14076:data <=32'h015AFFF0;14'd14077:data <=32'h015EFFA7;14'd14078:data <=32'h014DFF5A;
14'd14079:data <=32'h0127FF13;14'd14080:data <=32'h0085FF9F;14'd14081:data <=32'h008FFF81;
14'd14082:data <=32'h00A5FF65;14'd14083:data <=32'h00D9FF0D;14'd14084:data <=32'h006DFECD;
14'd14085:data <=32'h0033FECB;14'd14086:data <=32'hFFFFFED4;14'd14087:data <=32'hFFCFFEE6;
14'd14088:data <=32'hFFA5FF00;14'd14089:data <=32'hFF82FF22;14'd14090:data <=32'hFF6AFF49;
14'd14091:data <=32'hFF5FFF72;14'd14092:data <=32'hFF60FF96;14'd14093:data <=32'hFF68FFB4;
14'd14094:data <=32'hFF75FFCA;14'd14095:data <=32'hFF80FFD6;14'd14096:data <=32'hFF89FFDD;
14'd14097:data <=32'hFF8CFFE2;14'd14098:data <=32'hFF8DFFE9;14'd14099:data <=32'hFF8CFFF5;
14'd14100:data <=32'hFF8E0002;14'd14101:data <=32'hFF940010;14'd14102:data <=32'hFFA0001D;
14'd14103:data <=32'hFFAE0024;14'd14104:data <=32'hFFBD0025;14'd14105:data <=32'hFFC80022;
14'd14106:data <=32'hFFD0001C;14'd14107:data <=32'hFFD50015;14'd14108:data <=32'hFFD5000E;
14'd14109:data <=32'hFFD2000A;14'd14110:data <=32'hFFD10006;14'd14111:data <=32'hFFCD0004;
14'd14112:data <=32'hFFC70003;14'd14113:data <=32'hFFBF0003;14'd14114:data <=32'hFFB60006;
14'd14115:data <=32'hFFAB000E;14'd14116:data <=32'hFFA2001C;14'd14117:data <=32'hFF9E002D;
14'd14118:data <=32'hFF9F0043;14'd14119:data <=32'hFFAA0057;14'd14120:data <=32'hFFBC0068;
14'd14121:data <=32'hFFD20070;14'd14122:data <=32'hFFE9006E;14'd14123:data <=32'hFFFD0065;
14'd14124:data <=32'h00090056;14'd14125:data <=32'h000C0045;14'd14126:data <=32'h00070036;
14'd14127:data <=32'hFFFB002E;14'd14128:data <=32'hFFEC002D;14'd14129:data <=32'hFFDF0034;
14'd14130:data <=32'hFFD40042;14'd14131:data <=32'hFFCE0055;14'd14132:data <=32'hFFCD006C;
14'd14133:data <=32'hFFD30083;14'd14134:data <=32'hFFE1009E;14'd14135:data <=32'hFFF700B8;
14'd14136:data <=32'h001700CF;14'd14137:data <=32'h004100DF;14'd14138:data <=32'h007300E4;
14'd14139:data <=32'h00A900DA;14'd14140:data <=32'h00DE00BF;14'd14141:data <=32'h010A0094;
14'd14142:data <=32'h012A005D;14'd14143:data <=32'h01380020;14'd14144:data <=32'h010E004D;
14'd14145:data <=32'h0135001B;14'd14146:data <=32'h0143FFF7;14'd14147:data <=32'h010C000A;
14'd14148:data <=32'h00D2FFC0;14'd14149:data <=32'h00C6FFAC;14'd14150:data <=32'h00BBFF96;
14'd14151:data <=32'h00AEFF82;14'd14152:data <=32'h009FFF6D;14'd14153:data <=32'h008BFF5B;
14'd14154:data <=32'h0074FF4C;14'd14155:data <=32'h005DFF41;14'd14156:data <=32'h0045FF39;
14'd14157:data <=32'h002EFF32;14'd14158:data <=32'h0016FF2B;14'd14159:data <=32'hFFFAFF26;
14'd14160:data <=32'hFFD9FF24;14'd14161:data <=32'hFFB4FF2A;14'd14162:data <=32'hFF8EFF3A;
14'd14163:data <=32'hFF6CFF56;14'd14164:data <=32'hFF52FF7C;14'd14165:data <=32'hFF43FFAA;
14'd14166:data <=32'hFF45FFD7;14'd14167:data <=32'hFF520000;14'd14168:data <=32'hFF6B0021;
14'd14169:data <=32'hFF890036;14'd14170:data <=32'hFFA90040;14'd14171:data <=32'hFFC80041;
14'd14172:data <=32'hFFE20039;14'd14173:data <=32'hFFF6002C;14'd14174:data <=32'h0006001A;
14'd14175:data <=32'h000F0004;14'd14176:data <=32'h0011FFED;14'd14177:data <=32'h000AFFD6;
14'd14178:data <=32'hFFFBFFC1;14'd14179:data <=32'hFFE5FFB3;14'd14180:data <=32'hFFC9FFAD;
14'd14181:data <=32'hFFADFFB2;14'd14182:data <=32'hFF93FFC0;14'd14183:data <=32'hFF82FFD6;
14'd14184:data <=32'hFF78FFF0;14'd14185:data <=32'hFF78000A;14'd14186:data <=32'hFF7E001F;
14'd14187:data <=32'hFF89002F;14'd14188:data <=32'hFF930039;14'd14189:data <=32'hFF9A003D;
14'd14190:data <=32'hFF9F0042;14'd14191:data <=32'hFFA00049;14'd14192:data <=32'hFFA10050;
14'd14193:data <=32'hFFA2005D;14'd14194:data <=32'hFFA6006B;14'd14195:data <=32'hFFAE0079;
14'd14196:data <=32'hFFBA0087;14'd14197:data <=32'hFFC60093;14'd14198:data <=32'hFFD5009F;
14'd14199:data <=32'hFFE400AA;14'd14200:data <=32'hFFF800B2;14'd14201:data <=32'h001000BB;
14'd14202:data <=32'h002C00BF;14'd14203:data <=32'h004A00BD;14'd14204:data <=32'h006900B2;
14'd14205:data <=32'h0086009E;14'd14206:data <=32'h009B0083;14'd14207:data <=32'h00A70066;
14'd14208:data <=32'h007A0116;14'd14209:data <=32'h00C5010E;14'd14210:data <=32'h00F400E4;
14'd14211:data <=32'h008B0059;14'd14212:data <=32'h0056002C;14'd14213:data <=32'h00580038;
14'd14214:data <=32'h00620041;14'd14215:data <=32'h00750047;14'd14216:data <=32'h008B0043;
14'd14217:data <=32'h00A10036;14'd14218:data <=32'h00B50024;14'd14219:data <=32'h00C7000C;
14'd14220:data <=32'h00D5FFED;14'd14221:data <=32'h00DEFFCA;14'd14222:data <=32'h00DDFFA0;
14'd14223:data <=32'h00D3FF74;14'd14224:data <=32'h00BCFF47;14'd14225:data <=32'h0096FF1F;
14'd14226:data <=32'h0065FF02;14'd14227:data <=32'h002BFEF6;14'd14228:data <=32'hFFF1FEFB;
14'd14229:data <=32'hFFBBFF11;14'd14230:data <=32'hFF92FF34;14'd14231:data <=32'hFF76FF5E;
14'd14232:data <=32'hFF6AFF8B;14'd14233:data <=32'hFF68FFB4;14'd14234:data <=32'hFF72FFD8;
14'd14235:data <=32'hFF81FFF6;14'd14236:data <=32'hFF93000C;14'd14237:data <=32'hFFAB001D;
14'd14238:data <=32'hFFC30026;14'd14239:data <=32'hFFDE0029;14'd14240:data <=32'hFFF70024;
14'd14241:data <=32'h000D0017;14'd14242:data <=32'h001C0004;14'd14243:data <=32'h0024FFED;
14'd14244:data <=32'h0025FFD4;14'd14245:data <=32'h001BFFBE;14'd14246:data <=32'h000DFFAD;
14'd14247:data <=32'hFFFCFFA1;14'd14248:data <=32'hFFEBFF9A;14'd14249:data <=32'hFFD9FF96;
14'd14250:data <=32'hFFC9FF94;14'd14251:data <=32'hFFB7FF91;14'd14252:data <=32'hFFA2FF91;
14'd14253:data <=32'hFF89FF92;14'd14254:data <=32'hFF6EFF9A;14'd14255:data <=32'hFF4EFFAB;
14'd14256:data <=32'hFF32FFC6;14'd14257:data <=32'hFF1AFFEA;14'd14258:data <=32'hFF0E0016;
14'd14259:data <=32'hFF0C0044;14'd14260:data <=32'hFF180075;14'd14261:data <=32'hFF2E009F;
14'd14262:data <=32'hFF4C00C3;14'd14263:data <=32'hFF7100DE;14'd14264:data <=32'hFF9A00F4;
14'd14265:data <=32'hFFC600FF;14'd14266:data <=32'hFFF30101;14'd14267:data <=32'h002200FA;
14'd14268:data <=32'h004C00E7;14'd14269:data <=32'h007100C8;14'd14270:data <=32'h008900A1;
14'd14271:data <=32'h00930078;14'd14272:data <=32'hFFCA00D4;14'd14273:data <=32'hFFF200F5;
14'd14274:data <=32'h003100FA;14'd14275:data <=32'h0082006F;14'd14276:data <=32'h00440035;
14'd14277:data <=32'h0036003B;14'd14278:data <=32'h00300046;14'd14279:data <=32'h00340055;
14'd14280:data <=32'h003E005E;14'd14281:data <=32'h004D0065;14'd14282:data <=32'h005F0066;
14'd14283:data <=32'h00750064;14'd14284:data <=32'h008B005C;14'd14285:data <=32'h00A1004F;
14'd14286:data <=32'h00B70039;14'd14287:data <=32'h00C9001A;14'd14288:data <=32'h00D4FFF6;
14'd14289:data <=32'h00D2FFCB;14'd14290:data <=32'h00C4FFA4;14'd14291:data <=32'h00ABFF81;
14'd14292:data <=32'h008AFF69;14'd14293:data <=32'h0064FF5C;14'd14294:data <=32'h0043FF5C;
14'd14295:data <=32'h0025FF63;14'd14296:data <=32'h000EFF6D;14'd14297:data <=32'hFFFDFF79;
14'd14298:data <=32'hFFF0FF85;14'd14299:data <=32'hFFE5FF91;14'd14300:data <=32'hFFDBFF9B;
14'd14301:data <=32'hFFD1FFA8;14'd14302:data <=32'hFFC9FFB8;14'd14303:data <=32'hFFC7FFCA;
14'd14304:data <=32'hFFC9FFDB;14'd14305:data <=32'hFFD1FFEA;14'd14306:data <=32'hFFDCFFF7;
14'd14307:data <=32'hFFEAFFFC;14'd14308:data <=32'hFFF80000;14'd14309:data <=32'h0005FFFE;
14'd14310:data <=32'h0014FFFB;14'd14311:data <=32'h0021FFF3;14'd14312:data <=32'h002DFFE8;
14'd14313:data <=32'h0039FFD8;14'd14314:data <=32'h0043FFC2;14'd14315:data <=32'h0047FFA5;
14'd14316:data <=32'h0041FF83;14'd14317:data <=32'h002FFF5E;14'd14318:data <=32'h0010FF3D;
14'd14319:data <=32'hFFE4FF26;14'd14320:data <=32'hFFAEFF1B;14'd14321:data <=32'hFF75FF21;
14'd14322:data <=32'hFF3DFF39;14'd14323:data <=32'hFF0EFF5E;14'd14324:data <=32'hFEEAFF8F;
14'd14325:data <=32'hFED4FFC7;14'd14326:data <=32'hFECC0001;14'd14327:data <=32'hFED1003C;
14'd14328:data <=32'hFEE10073;14'd14329:data <=32'hFEFD00A4;14'd14330:data <=32'hFF2300CF;
14'd14331:data <=32'hFF5100EE;14'd14332:data <=32'hFF860102;14'd14333:data <=32'hFFBD0107;
14'd14334:data <=32'hFFEF00FC;14'd14335:data <=32'h001900E6;14'd14336:data <=32'hFFD00099;
14'd14337:data <=32'hFFDC00A6;14'd14338:data <=32'hFFEE00C1;14'd14339:data <=32'h001600F0;
14'd14340:data <=32'hFFFA00B6;14'd14341:data <=32'h000800B7;14'd14342:data <=32'h001A00BA;
14'd14343:data <=32'h003100BB;14'd14344:data <=32'h004A00B5;14'd14345:data <=32'h006200A8;
14'd14346:data <=32'h00770096;14'd14347:data <=32'h00880081;14'd14348:data <=32'h0092006B;
14'd14349:data <=32'h009B0054;14'd14350:data <=32'h009F003E;14'd14351:data <=32'h00A00028;
14'd14352:data <=32'h009F000F;14'd14353:data <=32'h0099FFF7;14'd14354:data <=32'h008CFFE2;
14'd14355:data <=32'h0079FFD1;14'd14356:data <=32'h0062FFC8;14'd14357:data <=32'h004DFFC7;
14'd14358:data <=32'h003CFFD0;14'd14359:data <=32'h0034FFDB;14'd14360:data <=32'h0033FFE7;
14'd14361:data <=32'h003AFFED;14'd14362:data <=32'h0045FFEE;14'd14363:data <=32'h004DFFE7;
14'd14364:data <=32'h0052FFDB;14'd14365:data <=32'h0050FFCC;14'd14366:data <=32'h0049FFBE;
14'd14367:data <=32'h003DFFB4;14'd14368:data <=32'h002FFFAF;14'd14369:data <=32'h0020FFAE;
14'd14370:data <=32'h0015FFB2;14'd14371:data <=32'h0009FFB7;14'd14372:data <=32'h0001FFC0;
14'd14373:data <=32'hFFFAFFCA;14'd14374:data <=32'hFFF9FFD6;14'd14375:data <=32'hFFFCFFE3;
14'd14376:data <=32'h0004FFF0;14'd14377:data <=32'h0014FFF8;14'd14378:data <=32'h0029FFFC;
14'd14379:data <=32'h003FFFF3;14'd14380:data <=32'h0056FFE1;14'd14381:data <=32'h0066FFC4;
14'd14382:data <=32'h006AFFA0;14'd14383:data <=32'h0061FF79;14'd14384:data <=32'h004BFF54;
14'd14385:data <=32'h0029FF39;14'd14386:data <=32'h0000FF27;14'd14387:data <=32'hFFD5FF21;
14'd14388:data <=32'hFFAAFF27;14'd14389:data <=32'hFF85FF35;14'd14390:data <=32'hFF62FF48;
14'd14391:data <=32'hFF45FF61;14'd14392:data <=32'hFF2CFF7E;14'd14393:data <=32'hFF18FF9F;
14'd14394:data <=32'hFF0AFFC3;14'd14395:data <=32'hFF04FFEA;14'd14396:data <=32'hFF070011;
14'd14397:data <=32'hFF100034;14'd14398:data <=32'hFF1F0052;14'd14399:data <=32'hFF31006A;
14'd14400:data <=32'hFF7700AF;14'd14401:data <=32'hFF8F00B9;14'd14402:data <=32'hFF9100B7;
14'd14403:data <=32'hFF200091;14'd14404:data <=32'hFEFE0086;14'd14405:data <=32'hFF0F00B7;
14'd14406:data <=32'hFF2E00E8;14'd14407:data <=32'hFF5A0113;14'd14408:data <=32'hFF920130;
14'd14409:data <=32'hFFD2013C;14'd14410:data <=32'h00100136;14'd14411:data <=32'h00480123;
14'd14412:data <=32'h00790104;14'd14413:data <=32'h009E00DD;14'd14414:data <=32'h00BA00B2;
14'd14415:data <=32'h00CA0083;14'd14416:data <=32'h00CF0053;14'd14417:data <=32'h00CA0025;
14'd14418:data <=32'h00B7FFFA;14'd14419:data <=32'h009BFFD8;14'd14420:data <=32'h0077FFC3;
14'd14421:data <=32'h0050FFBA;14'd14422:data <=32'h002CFFC0;14'd14423:data <=32'h0010FFD2;
14'd14424:data <=32'h0000FFEC;14'd14425:data <=32'hFFFD0006;14'd14426:data <=32'h0005001C;
14'd14427:data <=32'h0013002B;14'd14428:data <=32'h00260030;14'd14429:data <=32'h0036002F;
14'd14430:data <=32'h00430029;14'd14431:data <=32'h004C0020;14'd14432:data <=32'h00530016;
14'd14433:data <=32'h0058000D;14'd14434:data <=32'h005B0003;14'd14435:data <=32'h005DFFF8;
14'd14436:data <=32'h005CFFED;14'd14437:data <=32'h0058FFE4;14'd14438:data <=32'h0053FFDB;
14'd14439:data <=32'h004CFFD6;14'd14440:data <=32'h0046FFD4;14'd14441:data <=32'h0042FFD4;
14'd14442:data <=32'h0043FFD5;14'd14443:data <=32'h0047FFD4;14'd14444:data <=32'h004DFFCE;
14'd14445:data <=32'h0053FFC4;14'd14446:data <=32'h0055FFB5;14'd14447:data <=32'h0052FFA3;
14'd14448:data <=32'h0048FF92;14'd14449:data <=32'h0038FF84;14'd14450:data <=32'h0027FF7D;
14'd14451:data <=32'h0016FF7A;14'd14452:data <=32'h0007FF7E;14'd14453:data <=32'hFFFEFF82;
14'd14454:data <=32'hFFF9FF84;14'd14455:data <=32'hFFF6FF83;14'd14456:data <=32'hFFF1FF7C;
14'd14457:data <=32'hFFE8FF73;14'd14458:data <=32'hFFDBFF6A;14'd14459:data <=32'hFFCAFF62;
14'd14460:data <=32'hFFB3FF5C;14'd14461:data <=32'hFF9BFF59;14'd14462:data <=32'hFF7FFF5C;
14'd14463:data <=32'hFF62FF61;14'd14464:data <=32'hFF19FFFA;14'd14465:data <=32'hFF17000F;
14'd14466:data <=32'hFF260010;14'd14467:data <=32'hFF2EFF84;14'd14468:data <=32'hFEDAFF73;
14'd14469:data <=32'hFEB5FFAF;14'd14470:data <=32'hFEA0FFF4;14'd14471:data <=32'hFE9E003E;
14'd14472:data <=32'hFEB40087;14'd14473:data <=32'hFEDC00C7;14'd14474:data <=32'hFF0F00F7;
14'd14475:data <=32'hFF4C0118;14'd14476:data <=32'hFF880127;14'd14477:data <=32'hFFC4012A;
14'd14478:data <=32'hFFFC0121;14'd14479:data <=32'h0030010D;14'd14480:data <=32'h005C00EF;
14'd14481:data <=32'h007F00C9;14'd14482:data <=32'h0096009C;14'd14483:data <=32'h009F006D;
14'd14484:data <=32'h009A0041;14'd14485:data <=32'h0089001C;14'd14486:data <=32'h00710003;
14'd14487:data <=32'h0057FFF5;14'd14488:data <=32'h003EFFF1;14'd14489:data <=32'h002BFFF6;
14'd14490:data <=32'h001EFFFC;14'd14491:data <=32'h00160003;14'd14492:data <=32'h00120009;
14'd14493:data <=32'h000E000D;14'd14494:data <=32'h00090012;14'd14495:data <=32'h00040019;
14'd14496:data <=32'h00000024;14'd14497:data <=32'h00000032;14'd14498:data <=32'h00070040;
14'd14499:data <=32'h0011004D;14'd14500:data <=32'h00220057;14'd14501:data <=32'h0035005D;
14'd14502:data <=32'h004A005B;14'd14503:data <=32'h005E0055;14'd14504:data <=32'h0071004B;
14'd14505:data <=32'h0082003E;14'd14506:data <=32'h0091002C;14'd14507:data <=32'h009F0018;
14'd14508:data <=32'h00A9FFFF;14'd14509:data <=32'h00AFFFE1;14'd14510:data <=32'h00ABFFC2;
14'd14511:data <=32'h009FFFA2;14'd14512:data <=32'h008AFF87;14'd14513:data <=32'h006CFF72;
14'd14514:data <=32'h004BFF6A;14'd14515:data <=32'h002BFF6D;14'd14516:data <=32'h0011FF7A;
14'd14517:data <=32'h0002FF8E;14'd14518:data <=32'hFFFBFFA2;14'd14519:data <=32'h0001FFB3;
14'd14520:data <=32'h000DFFBC;14'd14521:data <=32'h001BFFBE;14'd14522:data <=32'h0027FFB5;
14'd14523:data <=32'h0031FFA6;14'd14524:data <=32'h0036FF92;14'd14525:data <=32'h0033FF7B;
14'd14526:data <=32'h002AFF61;14'd14527:data <=32'h0019FF47;14'd14528:data <=32'hFFCFFF57;
14'd14529:data <=32'hFFB8FF43;14'd14530:data <=32'hFFACFF45;14'd14531:data <=32'hFFDDFF52;
14'd14532:data <=32'hFF8AFF18;14'd14533:data <=32'hFF5BFF29;14'd14534:data <=32'hFF2FFF4A;
14'd14535:data <=32'hFF0DFF75;14'd14536:data <=32'hFEFBFFA8;14'd14537:data <=32'hFEF6FFDB;
14'd14538:data <=32'hFEFF0007;14'd14539:data <=32'hFF0E002D;14'd14540:data <=32'hFF21004C;
14'd14541:data <=32'hFF360067;14'd14542:data <=32'hFF4C007E;14'd14543:data <=32'hFF650090;
14'd14544:data <=32'hFF81009E;14'd14545:data <=32'hFF9E00A8;14'd14546:data <=32'hFFBC00AA;
14'd14547:data <=32'hFFD600A7;14'd14548:data <=32'hFFEE009E;14'd14549:data <=32'h00000092;
14'd14550:data <=32'h000E0087;14'd14551:data <=32'h0019007D;14'd14552:data <=32'h00230076;
14'd14553:data <=32'h002E006C;14'd14554:data <=32'h003B0060;14'd14555:data <=32'h0048004F;
14'd14556:data <=32'h004F003A;14'd14557:data <=32'h004F0023;14'd14558:data <=32'h0046000A;
14'd14559:data <=32'h0033FFF7;14'd14560:data <=32'h001AFFEB;14'd14561:data <=32'hFFFFFFEB;
14'd14562:data <=32'hFFE5FFF5;14'd14563:data <=32'hFFD20009;14'd14564:data <=32'hFFC70022;
14'd14565:data <=32'hFFC4003F;14'd14566:data <=32'hFFCC005A;14'd14567:data <=32'hFFDA0074;
14'd14568:data <=32'hFFEF0089;14'd14569:data <=32'h000B009A;14'd14570:data <=32'h002B00A3;
14'd14571:data <=32'h004F00A5;14'd14572:data <=32'h0075009D;14'd14573:data <=32'h0099008A;
14'd14574:data <=32'h00B8006D;14'd14575:data <=32'h00CD0047;14'd14576:data <=32'h00D7001D;
14'd14577:data <=32'h00D3FFF3;14'd14578:data <=32'h00C3FFCF;14'd14579:data <=32'h00AEFFB5;
14'd14580:data <=32'h0094FFA4;14'd14581:data <=32'h007DFF9E;14'd14582:data <=32'h006BFF9E;
14'd14583:data <=32'h0060FFA0;14'd14584:data <=32'h005BFFA2;14'd14585:data <=32'h0059FFA1;
14'd14586:data <=32'h0058FF9A;14'd14587:data <=32'h0056FF91;14'd14588:data <=32'h0052FF86;
14'd14589:data <=32'h004BFF7B;14'd14590:data <=32'h0042FF6E;14'd14591:data <=32'h0038FF60;
14'd14592:data <=32'h0075FFCA;14'd14593:data <=32'h008BFF98;14'd14594:data <=32'h007CFF6C;
14'd14595:data <=32'hFFFEFF60;14'd14596:data <=32'hFFBCFF2B;14'd14597:data <=32'hFF9BFF3D;
14'd14598:data <=32'hFF7FFF59;14'd14599:data <=32'hFF6DFF79;14'd14600:data <=32'hFF67FF9C;
14'd14601:data <=32'hFF6BFFBB;14'd14602:data <=32'hFF78FFD2;14'd14603:data <=32'hFF87FFDF;
14'd14604:data <=32'hFF94FFE4;14'd14605:data <=32'hFF9BFFE1;14'd14606:data <=32'hFF9CFFDE;
14'd14607:data <=32'hFF97FFDD;14'd14608:data <=32'hFF8EFFE0;14'd14609:data <=32'hFF86FFE7;
14'd14610:data <=32'hFF7DFFF1;14'd14611:data <=32'hFF76FFFF;14'd14612:data <=32'hFF71000E;
14'd14613:data <=32'hFF6E0020;14'd14614:data <=32'hFF6D0035;14'd14615:data <=32'hFF71004E;
14'd14616:data <=32'hFF7C0068;14'd14617:data <=32'hFF900081;14'd14618:data <=32'hFFAE0095;
14'd14619:data <=32'hFFD1009D;14'd14620:data <=32'hFFF6009B;14'd14621:data <=32'h0018008A;
14'd14622:data <=32'h00310070;14'd14623:data <=32'h003F0052;14'd14624:data <=32'h00400032;
14'd14625:data <=32'h00350017;14'd14626:data <=32'h00240002;14'd14627:data <=32'h000DFFF8;
14'd14628:data <=32'hFFF6FFF5;14'd14629:data <=32'hFFE1FFF9;14'd14630:data <=32'hFFD00005;
14'd14631:data <=32'hFFC10014;14'd14632:data <=32'hFFB70028;14'd14633:data <=32'hFFB2003E;
14'd14634:data <=32'hFFB30056;14'd14635:data <=32'hFFBC0071;14'd14636:data <=32'hFFCC0089;
14'd14637:data <=32'hFFE3009D;14'd14638:data <=32'hFFFF00A9;14'd14639:data <=32'h001F00AF;
14'd14640:data <=32'h003C00AC;14'd14641:data <=32'h005700A3;14'd14642:data <=32'h006D0096;
14'd14643:data <=32'h007F0089;14'd14644:data <=32'h008E007E;14'd14645:data <=32'h009F0073;
14'd14646:data <=32'h00B30067;14'd14647:data <=32'h00C90056;14'd14648:data <=32'h00E1003F;
14'd14649:data <=32'h00F5001D;14'd14650:data <=32'h0103FFF5;14'd14651:data <=32'h0107FFC9;
14'd14652:data <=32'h00FEFF99;14'd14653:data <=32'h00ECFF6D;14'd14654:data <=32'h00D0FF48;
14'd14655:data <=32'h00AEFF29;14'd14656:data <=32'h0050001D;14'd14657:data <=32'h0083000C;
14'd14658:data <=32'h00A9FFD5;14'd14659:data <=32'h0074FF16;14'd14660:data <=32'h001AFED5;
14'd14661:data <=32'hFFDFFEE5;14'd14662:data <=32'hFFADFF04;14'd14663:data <=32'hFF85FF2C;
14'd14664:data <=32'hFF6FFF5E;14'd14665:data <=32'hFF69FF8F;14'd14666:data <=32'hFF76FFBA;
14'd14667:data <=32'hFF8DFFD7;14'd14668:data <=32'hFFA6FFE8;14'd14669:data <=32'hFFC0FFEB;
14'd14670:data <=32'hFFD2FFE6;14'd14671:data <=32'hFFDCFFDA;14'd14672:data <=32'hFFDFFFCF;
14'd14673:data <=32'hFFDCFFC2;14'd14674:data <=32'hFFD5FFB9;14'd14675:data <=32'hFFC9FFB2;
14'd14676:data <=32'hFFBAFFAE;14'd14677:data <=32'hFFA9FFAF;14'd14678:data <=32'hFF94FFB5;
14'd14679:data <=32'hFF80FFC2;14'd14680:data <=32'hFF70FFD8;14'd14681:data <=32'hFF67FFF4;
14'd14682:data <=32'hFF670012;14'd14683:data <=32'hFF72002F;14'd14684:data <=32'hFF850045;
14'd14685:data <=32'hFF9D0054;14'd14686:data <=32'hFFB60057;14'd14687:data <=32'hFFCB0054;
14'd14688:data <=32'hFFDA004C;14'd14689:data <=32'hFFE30042;14'd14690:data <=32'hFFE80039;
14'd14691:data <=32'hFFEA0032;14'd14692:data <=32'hFFEB002E;14'd14693:data <=32'hFFEB002A;
14'd14694:data <=32'hFFED0026;14'd14695:data <=32'hFFED0021;14'd14696:data <=32'hFFEC001A;
14'd14697:data <=32'hFFE50015;14'd14698:data <=32'hFFDC0011;14'd14699:data <=32'hFFD10013;
14'd14700:data <=32'hFFC60017;14'd14701:data <=32'hFFBA0021;14'd14702:data <=32'hFFB1002D;
14'd14703:data <=32'hFFAC003D;14'd14704:data <=32'hFFA8004E;14'd14705:data <=32'hFFA60062;
14'd14706:data <=32'hFFA60079;14'd14707:data <=32'hFFAB0093;14'd14708:data <=32'hFFB600B3;
14'd14709:data <=32'hFFCB00D5;14'd14710:data <=32'hFFEE00F5;14'd14711:data <=32'h001D010E;
14'd14712:data <=32'h0059011B;14'd14713:data <=32'h00990116;14'd14714:data <=32'h00D800FE;
14'd14715:data <=32'h011200D4;14'd14716:data <=32'h013F009C;14'd14717:data <=32'h015C005B;
14'd14718:data <=32'h01680015;14'd14719:data <=32'h0165FFD0;14'd14720:data <=32'h0086001A;
14'd14721:data <=32'h00AA0012;14'd14722:data <=32'h00DE0003;14'd14723:data <=32'h0143FFA9;
14'd14724:data <=32'h00FFFF39;14'd14725:data <=32'h00CBFF18;14'd14726:data <=32'h0091FF06;
14'd14727:data <=32'h0059FF04;14'd14728:data <=32'h0027FF10;14'd14729:data <=32'h0001FF29;
14'd14730:data <=32'hFFE7FF44;14'd14731:data <=32'hFFDAFF5F;14'd14732:data <=32'hFFD7FF75;
14'd14733:data <=32'hFFD5FF83;14'd14734:data <=32'hFFD3FF8C;14'd14735:data <=32'hFFD1FF93;
14'd14736:data <=32'hFFCAFF9A;14'd14737:data <=32'hFFC5FFA2;14'd14738:data <=32'hFFC1FFAC;
14'd14739:data <=32'hFFBFFFB4;14'd14740:data <=32'hFFBFFFBC;14'd14741:data <=32'hFFC0FFC2;
14'd14742:data <=32'hFFBFFFC6;14'd14743:data <=32'hFFBCFFCA;14'd14744:data <=32'hFFB9FFCF;
14'd14745:data <=32'hFFB6FFD7;14'd14746:data <=32'hFFB6FFDF;14'd14747:data <=32'hFFB9FFE8;
14'd14748:data <=32'hFFBEFFEE;14'd14749:data <=32'hFFC7FFF0;14'd14750:data <=32'hFFCDFFED;
14'd14751:data <=32'hFFCDFFE7;14'd14752:data <=32'hFFC9FFDF;14'd14753:data <=32'hFFBEFFDB;
14'd14754:data <=32'hFFB1FFDD;14'd14755:data <=32'hFFA4FFE6;14'd14756:data <=32'hFF9AFFF6;
14'd14757:data <=32'hFF980007;14'd14758:data <=32'hFF9B0019;14'd14759:data <=32'hFFA60027;
14'd14760:data <=32'hFFB30031;14'd14761:data <=32'hFFC20033;14'd14762:data <=32'hFFCF0030;
14'd14763:data <=32'hFFD8002A;14'd14764:data <=32'hFFDB0020;14'd14765:data <=32'hFFDC0017;
14'd14766:data <=32'hFFD8000D;14'd14767:data <=32'hFFCF0006;14'd14768:data <=32'hFFC10001;
14'd14769:data <=32'hFFAF0000;14'd14770:data <=32'hFF990005;14'd14771:data <=32'hFF800013;
14'd14772:data <=32'hFF6A002F;14'd14773:data <=32'hFF5B0055;14'd14774:data <=32'hFF560084;
14'd14775:data <=32'hFF6200B7;14'd14776:data <=32'hFF8000E8;14'd14777:data <=32'hFFAD0111;
14'd14778:data <=32'hFFE6012B;14'd14779:data <=32'h00240134;14'd14780:data <=32'h0062012D;
14'd14781:data <=32'h009B0118;14'd14782:data <=32'h00CC00F7;14'd14783:data <=32'h00F400CE;
14'd14784:data <=32'h00AD00CB;14'd14785:data <=32'h00E600BE;14'd14786:data <=32'h010C00B3;
14'd14787:data <=32'h00F400B8;14'd14788:data <=32'h00E80054;14'd14789:data <=32'h00EC0030;
14'd14790:data <=32'h00E80010;14'd14791:data <=32'h00E1FFF1;14'd14792:data <=32'h00D6FFDA;
14'd14793:data <=32'h00CBFFC8;14'd14794:data <=32'h00C3FFB6;14'd14795:data <=32'h00BDFFA3;
14'd14796:data <=32'h00B7FF8B;14'd14797:data <=32'h00AAFF6F;14'd14798:data <=32'h0096FF53;
14'd14799:data <=32'h0078FF39;14'd14800:data <=32'h0052FF29;14'd14801:data <=32'h0026FF22;
14'd14802:data <=32'hFFFDFF29;14'd14803:data <=32'hFFD7FF39;14'd14804:data <=32'hFFB9FF51;
14'd14805:data <=32'hFFA3FF6E;14'd14806:data <=32'hFF96FF8B;14'd14807:data <=32'hFF90FFA9;
14'd14808:data <=32'hFF90FFC7;14'd14809:data <=32'hFF98FFE3;14'd14810:data <=32'hFFA6FFFB;
14'd14811:data <=32'hFFBB000D;14'd14812:data <=32'hFFD50017;14'd14813:data <=32'hFFF10018;
14'd14814:data <=32'h000B000D;14'd14815:data <=32'h001DFFF9;14'd14816:data <=32'h0025FFDE;
14'd14817:data <=32'h0021FFC1;14'd14818:data <=32'h0014FFAB;14'd14819:data <=32'hFFFEFF9A;
14'd14820:data <=32'hFFE4FF96;14'd14821:data <=32'hFFCBFF97;14'd14822:data <=32'hFFB7FFA1;
14'd14823:data <=32'hFFA8FFB0;14'd14824:data <=32'hFFA0FFBF;14'd14825:data <=32'hFF9CFFCD;
14'd14826:data <=32'hFF99FFD8;14'd14827:data <=32'hFF99FFE3;14'd14828:data <=32'hFF97FFEB;
14'd14829:data <=32'hFF98FFF2;14'd14830:data <=32'hFF98FFF9;14'd14831:data <=32'hFF98FFFE;
14'd14832:data <=32'hFF970002;14'd14833:data <=32'hFF960005;14'd14834:data <=32'hFF900009;
14'd14835:data <=32'hFF86000E;14'd14836:data <=32'hFF7A0017;14'd14837:data <=32'hFF6D0028;
14'd14838:data <=32'hFF640041;14'd14839:data <=32'hFF640060;14'd14840:data <=32'hFF6D0080;
14'd14841:data <=32'hFF7F00A0;14'd14842:data <=32'hFF9B00B8;14'd14843:data <=32'hFFBB00C6;
14'd14844:data <=32'hFFDA00CC;14'd14845:data <=32'hFFF800C8;14'd14846:data <=32'h001000C4;
14'd14847:data <=32'h002400BC;14'd14848:data <=32'hFFD1013B;14'd14849:data <=32'h0014015F;
14'd14850:data <=32'h00510157;14'd14851:data <=32'h002400C6;14'd14852:data <=32'h00170088;
14'd14853:data <=32'h001F0091;14'd14854:data <=32'h002D0099;14'd14855:data <=32'h003F00A0;
14'd14856:data <=32'h005400A7;14'd14857:data <=32'h007000AC;14'd14858:data <=32'h009400A9;
14'd14859:data <=32'h00BB009C;14'd14860:data <=32'h00E30082;14'd14861:data <=32'h01060058;
14'd14862:data <=32'h011C0023;14'd14863:data <=32'h0123FFE6;14'd14864:data <=32'h0116FFAA;
14'd14865:data <=32'h00F9FF75;14'd14866:data <=32'h00D0FF4B;14'd14867:data <=32'h009FFF2F;
14'd14868:data <=32'h006DFF21;14'd14869:data <=32'h003BFF20;14'd14870:data <=32'h000EFF29;
14'd14871:data <=32'hFFE6FF3B;14'd14872:data <=32'hFFC5FF56;14'd14873:data <=32'hFFACFF76;
14'd14874:data <=32'hFF9CFF9B;14'd14875:data <=32'hFF98FFC2;14'd14876:data <=32'hFFA1FFE7;
14'd14877:data <=32'hFFB50005;14'd14878:data <=32'hFFD00018;14'd14879:data <=32'hFFEF001F;
14'd14880:data <=32'h000B001C;14'd14881:data <=32'h0022000F;14'd14882:data <=32'h0031FFFD;
14'd14883:data <=32'h0039FFEA;14'd14884:data <=32'h003BFFD6;14'd14885:data <=32'h0038FFC6;
14'd14886:data <=32'h0034FFB8;14'd14887:data <=32'h002EFFAB;14'd14888:data <=32'h0029FF9D;
14'd14889:data <=32'h0020FF8E;14'd14890:data <=32'h0013FF7E;14'd14891:data <=32'h0002FF6E;
14'd14892:data <=32'hFFEAFF62;14'd14893:data <=32'hFFCDFF5C;14'd14894:data <=32'hFFADFF5B;
14'd14895:data <=32'hFF8FFF63;14'd14896:data <=32'hFF71FF71;14'd14897:data <=32'hFF57FF85;
14'd14898:data <=32'hFF41FF9E;14'd14899:data <=32'hFF2DFFBA;14'd14900:data <=32'hFF1FFFDA;
14'd14901:data <=32'hFF16FFFE;14'd14902:data <=32'hFF140027;14'd14903:data <=32'hFF1D0051;
14'd14904:data <=32'hFF30007A;14'd14905:data <=32'hFF4F009D;14'd14906:data <=32'hFF7700B5;
14'd14907:data <=32'hFFA200BE;14'd14908:data <=32'hFFCA00BA;14'd14909:data <=32'hFFEA00AA;
14'd14910:data <=32'h00000092;14'd14911:data <=32'h000A007C;14'd14912:data <=32'hFF3A0095;
14'd14913:data <=32'hFF4700D0;14'd14914:data <=32'hFF7C00F9;14'd14915:data <=32'hFFFD0093;
14'd14916:data <=32'hFFE3004F;14'd14917:data <=32'hFFD80055;14'd14918:data <=32'hFFD00060;
14'd14919:data <=32'hFFCF0072;14'd14920:data <=32'hFFD00087;14'd14921:data <=32'hFFDA00A1;
14'd14922:data <=32'hFFF000BA;14'd14923:data <=32'h001100CF;14'd14924:data <=32'h003D00D9;
14'd14925:data <=32'h006C00D4;14'd14926:data <=32'h009A00C1;14'd14927:data <=32'h00C1009F;
14'd14928:data <=32'h00DB0074;14'd14929:data <=32'h00E80045;14'd14930:data <=32'h00E70017;
14'd14931:data <=32'h00DBFFEF;14'd14932:data <=32'h00CAFFCE;14'd14933:data <=32'h00B5FFB4;
14'd14934:data <=32'h009EFF9E;14'd14935:data <=32'h0084FF8E;14'd14936:data <=32'h0068FF82;
14'd14937:data <=32'h004CFF7D;14'd14938:data <=32'h002FFF7F;14'd14939:data <=32'h0015FF88;
14'd14940:data <=32'h0000FF97;14'd14941:data <=32'hFFF1FFAA;14'd14942:data <=32'hFFEBFFBD;
14'd14943:data <=32'hFFEAFFCF;14'd14944:data <=32'hFFEDFFDD;14'd14945:data <=32'hFFF2FFE9;
14'd14946:data <=32'hFFF7FFF1;14'd14947:data <=32'hFFFCFFF9;14'd14948:data <=32'h00040002;
14'd14949:data <=32'h000F000C;14'd14950:data <=32'h001E0013;14'd14951:data <=32'h00340017;
14'd14952:data <=32'h004E0011;14'd14953:data <=32'h00690003;14'd14954:data <=32'h0080FFE9;
14'd14955:data <=32'h008EFFC4;14'd14956:data <=32'h0092FF9B;14'd14957:data <=32'h0088FF70;
14'd14958:data <=32'h0070FF47;14'd14959:data <=32'h004EFF24;14'd14960:data <=32'h0025FF0B;
14'd14961:data <=32'hFFF5FEFD;14'd14962:data <=32'hFFC2FEF8;14'd14963:data <=32'hFF8DFEFE;
14'd14964:data <=32'hFF5AFF11;14'd14965:data <=32'hFF29FF31;14'd14966:data <=32'hFF02FF5D;
14'd14967:data <=32'hFEE4FF92;14'd14968:data <=32'hFED8FFCE;14'd14969:data <=32'hFEDC000A;
14'd14970:data <=32'hFEF10042;14'd14971:data <=32'hFF12006E;14'd14972:data <=32'hFF3D008B;
14'd14973:data <=32'hFF670098;14'd14974:data <=32'hFF8D0098;14'd14975:data <=32'hFFAA008F;
14'd14976:data <=32'hFF7A0031;14'd14977:data <=32'hFF6D0045;14'd14978:data <=32'hFF6A006F;
14'd14979:data <=32'hFF9200B4;14'd14980:data <=32'hFF8E0079;14'd14981:data <=32'hFF9A0082;
14'd14982:data <=32'hFFA6008B;14'd14983:data <=32'hFFB30093;14'd14984:data <=32'hFFBF009A;
14'd14985:data <=32'hFFCC00A2;14'd14986:data <=32'hFFDE00AB;14'd14987:data <=32'hFFF300B4;
14'd14988:data <=32'h000E00B8;14'd14989:data <=32'h002B00B4;14'd14990:data <=32'h004800A9;
14'd14991:data <=32'h00610092;14'd14992:data <=32'h00700078;14'd14993:data <=32'h0076005C;
14'd14994:data <=32'h00730045;14'd14995:data <=32'h006B0033;14'd14996:data <=32'h0061002A;
14'd14997:data <=32'h00590025;14'd14998:data <=32'h00560024;14'd14999:data <=32'h00580022;
14'd15000:data <=32'h005B001D;14'd15001:data <=32'h005E0017;14'd15002:data <=32'h0060000E;
14'd15003:data <=32'h00600004;14'd15004:data <=32'h005EFFFC;14'd15005:data <=32'h005CFFF4;
14'd15006:data <=32'h0059FFEA;14'd15007:data <=32'h0055FFE0;14'd15008:data <=32'h004EFFD6;
14'd15009:data <=32'h0044FFCE;14'd15010:data <=32'h0036FFC6;14'd15011:data <=32'h0023FFC4;
14'd15012:data <=32'h0011FFCB;14'd15013:data <=32'h0002FFD9;14'd15014:data <=32'hFFFAFFEF;
14'd15015:data <=32'hFFFC0008;14'd15016:data <=32'h0009001F;14'd15017:data <=32'h00210030;
14'd15018:data <=32'h00410036;14'd15019:data <=32'h00630031;14'd15020:data <=32'h0081001E;
14'd15021:data <=32'h009A0002;14'd15022:data <=32'h00A9FFDE;14'd15023:data <=32'h00AEFFB8;
14'd15024:data <=32'h00A9FF90;14'd15025:data <=32'h009CFF6A;14'd15026:data <=32'h0087FF47;
14'd15027:data <=32'h0068FF28;14'd15028:data <=32'h0043FF0F;14'd15029:data <=32'h0017FEFE;
14'd15030:data <=32'hFFE8FEF8;14'd15031:data <=32'hFFB7FEFF;14'd15032:data <=32'hFF8AFF11;
14'd15033:data <=32'hFF66FF2D;14'd15034:data <=32'hFF4AFF4F;14'd15035:data <=32'hFF3BFF72;
14'd15036:data <=32'hFF34FF91;14'd15037:data <=32'hFF32FFAC;14'd15038:data <=32'hFF31FFC1;
14'd15039:data <=32'hFF2EFFD4;14'd15040:data <=32'hFF5F002C;14'd15041:data <=32'hFF630034;
14'd15042:data <=32'hFF580034;14'd15043:data <=32'hFEF10000;14'd15044:data <=32'hFED9FFEE;
14'd15045:data <=32'hFED70022;14'd15046:data <=32'hFEE20056;14'd15047:data <=32'hFEF80087;
14'd15048:data <=32'hFF1700AF;14'd15049:data <=32'hFF3C00CF;14'd15050:data <=32'hFF6700EB;
14'd15051:data <=32'hFF9700FC;14'd15052:data <=32'hFFCB0103;14'd15053:data <=32'hFFFF00FC;
14'd15054:data <=32'h003100E8;14'd15055:data <=32'h005900C6;14'd15056:data <=32'h0073009B;
14'd15057:data <=32'h007E006E;14'd15058:data <=32'h00780043;14'd15059:data <=32'h00660022;
14'd15060:data <=32'h004C000D;14'd15061:data <=32'h00320004;14'd15062:data <=32'h001B0006;
14'd15063:data <=32'h000B0010;14'd15064:data <=32'h0002001E;14'd15065:data <=32'hFFFF002B;
14'd15066:data <=32'h00010036;14'd15067:data <=32'h00070041;14'd15068:data <=32'h0010004A;
14'd15069:data <=32'h001C0050;14'd15070:data <=32'h002B0053;14'd15071:data <=32'h003C0051;
14'd15072:data <=32'h004B0049;14'd15073:data <=32'h0058003A;14'd15074:data <=32'h005F002A;
14'd15075:data <=32'h005D0018;14'd15076:data <=32'h00570008;14'd15077:data <=32'h004BFFFF;
14'd15078:data <=32'h0040FFFD;14'd15079:data <=32'h00350001;14'd15080:data <=32'h0032000A;
14'd15081:data <=32'h00350015;14'd15082:data <=32'h003E001C;14'd15083:data <=32'h004C001F;
14'd15084:data <=32'h00590019;14'd15085:data <=32'h0066000F;14'd15086:data <=32'h006E0004;
14'd15087:data <=32'h0073FFF6;14'd15088:data <=32'h0075FFE9;14'd15089:data <=32'h0077FFDC;
14'd15090:data <=32'h0077FFD1;14'd15091:data <=32'h0078FFC5;14'd15092:data <=32'h0078FFB5;
14'd15093:data <=32'h0076FFA5;14'd15094:data <=32'h0070FF94;14'd15095:data <=32'h0068FF82;
14'd15096:data <=32'h005EFF73;14'd15097:data <=32'h0051FF66;14'd15098:data <=32'h0045FF5A;
14'd15099:data <=32'h003AFF4C;14'd15100:data <=32'h002DFF3A;14'd15101:data <=32'h001AFF27;
14'd15102:data <=32'h0000FF10;14'd15103:data <=32'hFFDBFEFE;14'd15104:data <=32'hFF5EFF8A;
14'd15105:data <=32'hFF52FF94;14'd15106:data <=32'hFF57FF91;14'd15107:data <=32'hFF7EFF0A;
14'd15108:data <=32'hFF34FEDF;14'd15109:data <=32'hFEFCFF0A;14'd15110:data <=32'hFECFFF42;
14'd15111:data <=32'hFEB2FF83;14'd15112:data <=32'hFEA5FFC7;14'd15113:data <=32'hFEA60008;
14'd15114:data <=32'hFEB40049;14'd15115:data <=32'hFED10084;14'd15116:data <=32'hFEFC00B8;
14'd15117:data <=32'hFF3100DE;14'd15118:data <=32'hFF6F00F5;14'd15119:data <=32'hFFAE00F8;
14'd15120:data <=32'hFFE600E9;14'd15121:data <=32'h001400CE;14'd15122:data <=32'h003200A9;
14'd15123:data <=32'h00410083;14'd15124:data <=32'h00450060;14'd15125:data <=32'h003F0046;
14'd15126:data <=32'h00340032;14'd15127:data <=32'h00290026;14'd15128:data <=32'h001F001D;
14'd15129:data <=32'h00140017;14'd15130:data <=32'h000C0014;14'd15131:data <=32'h00000013;
14'd15132:data <=32'hFFF50015;14'd15133:data <=32'hFFED001B;14'd15134:data <=32'hFFE50026;
14'd15135:data <=32'hFFE40032;14'd15136:data <=32'hFFE6003F;14'd15137:data <=32'hFFEB0048;
14'd15138:data <=32'hFFF40051;14'd15139:data <=32'hFFFC0057;14'd15140:data <=32'h0004005A;
14'd15141:data <=32'h000B005F;14'd15142:data <=32'h00130065;14'd15143:data <=32'h001E006B;
14'd15144:data <=32'h002F0071;14'd15145:data <=32'h00420074;14'd15146:data <=32'h005A0071;
14'd15147:data <=32'h00720064;14'd15148:data <=32'h00870052;14'd15149:data <=32'h00950037;
14'd15150:data <=32'h009A001B;14'd15151:data <=32'h0095FFFF;14'd15152:data <=32'h0089FFE9;
14'd15153:data <=32'h0078FFDA;14'd15154:data <=32'h0066FFD3;14'd15155:data <=32'h0058FFD4;
14'd15156:data <=32'h004CFFD7;14'd15157:data <=32'h0048FFDF;14'd15158:data <=32'h0047FFE6;
14'd15159:data <=32'h004AFFEC;14'd15160:data <=32'h0053FFF1;14'd15161:data <=32'h0060FFF3;
14'd15162:data <=32'h0072FFF1;14'd15163:data <=32'h0087FFE6;14'd15164:data <=32'h009EFFD1;
14'd15165:data <=32'h00B1FFB1;14'd15166:data <=32'h00BBFF84;14'd15167:data <=32'h00B7FF50;
14'd15168:data <=32'h0046FF4E;14'd15169:data <=32'h0038FF2B;14'd15170:data <=32'h002BFF23;
14'd15171:data <=32'h005EFF32;14'd15172:data <=32'h0024FEDB;14'd15173:data <=32'hFFECFED7;
14'd15174:data <=32'hFFB8FEE1;14'd15175:data <=32'hFF86FEF6;14'd15176:data <=32'hFF5EFF13;
14'd15177:data <=32'hFF3CFF34;14'd15178:data <=32'hFF20FF5B;14'd15179:data <=32'hFF0DFF87;
14'd15180:data <=32'hFF03FFB5;14'd15181:data <=32'hFF05FFE4;14'd15182:data <=32'hFF12000F;
14'd15183:data <=32'hFF290032;14'd15184:data <=32'hFF44004B;14'd15185:data <=32'hFF60005A;
14'd15186:data <=32'hFF780062;14'd15187:data <=32'hFF8C0065;14'd15188:data <=32'hFF9C0068;
14'd15189:data <=32'hFFA8006B;14'd15190:data <=32'hFFB70071;14'd15191:data <=32'hFFCA0075;
14'd15192:data <=32'hFFDE0077;14'd15193:data <=32'hFFF40073;14'd15194:data <=32'h00080067;
14'd15195:data <=32'h00180055;14'd15196:data <=32'h00220040;14'd15197:data <=32'h0021002A;
14'd15198:data <=32'h001B0017;14'd15199:data <=32'h00100007;14'd15200:data <=32'hFFFFFFFE;
14'd15201:data <=32'hFFEFFFF8;14'd15202:data <=32'hFFDDFFF9;14'd15203:data <=32'hFFCCFFFE;
14'd15204:data <=32'hFFB9000A;14'd15205:data <=32'hFFAA001C;14'd15206:data <=32'hFF9E0034;
14'd15207:data <=32'hFF9B0053;14'd15208:data <=32'hFFA10074;14'd15209:data <=32'hFFB30094;
14'd15210:data <=32'hFFD100AF;14'd15211:data <=32'hFFF600C0;14'd15212:data <=32'h002000C4;
14'd15213:data <=32'h004900BB;14'd15214:data <=32'h006B00A6;14'd15215:data <=32'h0083008A;
14'd15216:data <=32'h0091006C;14'd15217:data <=32'h0096004E;14'd15218:data <=32'h00930035;
14'd15219:data <=32'h008C0023;14'd15220:data <=32'h00840016;14'd15221:data <=32'h007D000D;
14'd15222:data <=32'h00770006;14'd15223:data <=32'h00710001;14'd15224:data <=32'h006D0001;
14'd15225:data <=32'h006D0002;14'd15226:data <=32'h00710005;14'd15227:data <=32'h007B0005;
14'd15228:data <=32'h008B0000;14'd15229:data <=32'h009EFFF5;14'd15230:data <=32'h00B1FFDF;
14'd15231:data <=32'h00BDFFBE;14'd15232:data <=32'h00B7001A;14'd15233:data <=32'h00E2FFEC;
14'd15234:data <=32'h00E5FFBA;14'd15235:data <=32'h007BFF8D;14'd15236:data <=32'h0055FF3D;
14'd15237:data <=32'h0033FF3D;14'd15238:data <=32'h0016FF43;14'd15239:data <=32'h0000FF50;
14'd15240:data <=32'hFFF0FF5C;14'd15241:data <=32'hFFE5FF66;14'd15242:data <=32'hFFDCFF6E;
14'd15243:data <=32'hFFD2FF74;14'd15244:data <=32'hFFC9FF7B;14'd15245:data <=32'hFFC0FF82;
14'd15246:data <=32'hFFBAFF89;14'd15247:data <=32'hFFB3FF8E;14'd15248:data <=32'hFFACFF92;
14'd15249:data <=32'hFFA2FF93;14'd15250:data <=32'hFF94FF95;14'd15251:data <=32'hFF81FF9A;
14'd15252:data <=32'hFF6BFFA7;14'd15253:data <=32'hFF56FFBD;14'd15254:data <=32'hFF46FFDE;
14'd15255:data <=32'hFF420004;14'd15256:data <=32'hFF49002A;14'd15257:data <=32'hFF5D004C;
14'd15258:data <=32'hFF7A0066;14'd15259:data <=32'hFF9D0076;14'd15260:data <=32'hFFBF0077;
14'd15261:data <=32'hFFDE0071;14'd15262:data <=32'hFFF80062;14'd15263:data <=32'h000C004E;
14'd15264:data <=32'h00170038;14'd15265:data <=32'h001A0021;14'd15266:data <=32'h00180008;
14'd15267:data <=32'h000DFFF2;14'd15268:data <=32'hFFFCFFE1;14'd15269:data <=32'hFFE3FFD6;
14'd15270:data <=32'hFFC7FFD3;14'd15271:data <=32'hFFA9FFDC;14'd15272:data <=32'hFF90FFEF;
14'd15273:data <=32'hFF7D000A;14'd15274:data <=32'hFF74002C;14'd15275:data <=32'hFF78004E;
14'd15276:data <=32'hFF84006C;14'd15277:data <=32'hFF970085;14'd15278:data <=32'hFFAD0096;
14'd15279:data <=32'hFFC300A0;14'd15280:data <=32'hFFD700A6;14'd15281:data <=32'hFFE900AC;
14'd15282:data <=32'hFFFB00B2;14'd15283:data <=32'h000F00B8;14'd15284:data <=32'h002600BD;
14'd15285:data <=32'h004000BF;14'd15286:data <=32'h005D00BC;14'd15287:data <=32'h007A00B3;
14'd15288:data <=32'h009700A4;14'd15289:data <=32'h00AF0090;14'd15290:data <=32'h00C50079;
14'd15291:data <=32'h00D7005F;14'd15292:data <=32'h00E70042;14'd15293:data <=32'h00F40021;
14'd15294:data <=32'h00FCFFFA;14'd15295:data <=32'h00FCFFD0;14'd15296:data <=32'h004D0080;
14'd15297:data <=32'h008C0081;14'd15298:data <=32'h00C70059;14'd15299:data <=32'h00CDFF8E;
14'd15300:data <=32'h0099FF34;14'd15301:data <=32'h0065FF2E;14'd15302:data <=32'h0037FF3B;
14'd15303:data <=32'h0011FF52;14'd15304:data <=32'hFFFBFF6C;14'd15305:data <=32'hFFF0FF87;
14'd15306:data <=32'hFFEFFF9E;14'd15307:data <=32'hFFF4FFAF;14'd15308:data <=32'hFFFBFFBB;
14'd15309:data <=32'h0005FFC2;14'd15310:data <=32'h0011FFC3;14'd15311:data <=32'h001CFFBE;
14'd15312:data <=32'h0026FFB2;14'd15313:data <=32'h0029FF9F;14'd15314:data <=32'h0025FF89;
14'd15315:data <=32'h0015FF72;14'd15316:data <=32'hFFFAFF60;14'd15317:data <=32'hFFD8FF58;
14'd15318:data <=32'hFFB3FF5E;14'd15319:data <=32'hFF92FF6F;14'd15320:data <=32'hFF77FF8A;
14'd15321:data <=32'hFF69FFAC;14'd15322:data <=32'hFF65FFCD;14'd15323:data <=32'hFF6AFFEB;
14'd15324:data <=32'hFF770003;14'd15325:data <=32'hFF860016;14'd15326:data <=32'hFF970023;
14'd15327:data <=32'hFFA7002B;14'd15328:data <=32'hFFB80030;14'd15329:data <=32'hFFC90030;
14'd15330:data <=32'hFFD9002E;14'd15331:data <=32'hFFE70026;14'd15332:data <=32'hFFF1001A;
14'd15333:data <=32'hFFF6000B;14'd15334:data <=32'hFFF5FFFC;14'd15335:data <=32'hFFEEFFEE;
14'd15336:data <=32'hFFE2FFE4;14'd15337:data <=32'hFFD4FFDF;14'd15338:data <=32'hFFC6FFDF;
14'd15339:data <=32'hFFB9FFE2;14'd15340:data <=32'hFFAEFFE6;14'd15341:data <=32'hFFA3FFEB;
14'd15342:data <=32'hFF96FFF0;14'd15343:data <=32'hFF85FFF6;14'd15344:data <=32'hFF740002;
14'd15345:data <=32'hFF5F0016;14'd15346:data <=32'hFF4D0032;14'd15347:data <=32'hFF400059;
14'd15348:data <=32'hFF400086;14'd15349:data <=32'hFF4C00B9;14'd15350:data <=32'hFF6900E7;
14'd15351:data <=32'hFF90010F;14'd15352:data <=32'hFFC3012D;14'd15353:data <=32'hFFFC013E;
14'd15354:data <=32'h00380142;14'd15355:data <=32'h0075013A;14'd15356:data <=32'h00B00125;
14'd15357:data <=32'h00E80103;14'd15358:data <=32'h011800D4;14'd15359:data <=32'h013D0098;
14'd15360:data <=32'h0046007D;14'd15361:data <=32'h006F008B;14'd15362:data <=32'h00AC0093;
14'd15363:data <=32'h01370053;14'd15364:data <=32'h0122FFD4;14'd15365:data <=32'h00FEFFA8;
14'd15366:data <=32'h00D5FF8C;14'd15367:data <=32'h00ABFF7E;14'd15368:data <=32'h0088FF7B;
14'd15369:data <=32'h006CFF7D;14'd15370:data <=32'h0056FF84;14'd15371:data <=32'h0046FF8A;
14'd15372:data <=32'h0038FF92;14'd15373:data <=32'h002DFF9A;14'd15374:data <=32'h0026FFA1;
14'd15375:data <=32'h0024FFAA;14'd15376:data <=32'h0025FFAF;14'd15377:data <=32'h0028FFAF;
14'd15378:data <=32'h0029FFA9;14'd15379:data <=32'h0027FFA0;14'd15380:data <=32'h0020FF95;
14'd15381:data <=32'h0012FF8C;14'd15382:data <=32'h0001FF8B;14'd15383:data <=32'hFFEFFF8E;
14'd15384:data <=32'hFFDFFF98;14'd15385:data <=32'hFFD7FFA5;14'd15386:data <=32'hFFD3FFB2;
14'd15387:data <=32'hFFD5FFBB;14'd15388:data <=32'hFFD8FFC0;14'd15389:data <=32'hFFDBFFC1;
14'd15390:data <=32'hFFD9FFC0;14'd15391:data <=32'hFFD5FFBD;14'd15392:data <=32'hFFCDFFBE;
14'd15393:data <=32'hFFC4FFC2;14'd15394:data <=32'hFFBCFFCA;14'd15395:data <=32'hFFB9FFD3;
14'd15396:data <=32'hFFB7FFDC;14'd15397:data <=32'hFFB8FFE6;14'd15398:data <=32'hFFBBFFED;
14'd15399:data <=32'hFFBFFFF3;14'd15400:data <=32'hFFC4FFF8;14'd15401:data <=32'hFFCAFFFB;
14'd15402:data <=32'hFFD1FFFD;14'd15403:data <=32'hFFDAFFFB;14'd15404:data <=32'hFFE3FFF5;
14'd15405:data <=32'hFFEAFFE8;14'd15406:data <=32'hFFEAFFD5;14'd15407:data <=32'hFFE1FFC0;
14'd15408:data <=32'hFFCDFFAA;14'd15409:data <=32'hFFAFFF9D;14'd15410:data <=32'hFF86FF9B;
14'd15411:data <=32'hFF5BFFA7;14'd15412:data <=32'hFF32FFC3;14'd15413:data <=32'hFF12FFEC;
14'd15414:data <=32'hFEFF001F;14'd15415:data <=32'hFEF90059;14'd15416:data <=32'hFF030092;
14'd15417:data <=32'hFF1B00C8;14'd15418:data <=32'hFF3E00F8;14'd15419:data <=32'hFF6A011F;
14'd15420:data <=32'hFFA1013D;14'd15421:data <=32'hFFDC014F;14'd15422:data <=32'h001E0153;
14'd15423:data <=32'h005E0147;14'd15424:data <=32'h00220102;14'd15425:data <=32'h00580111;
14'd15426:data <=32'h007E011B;14'd15427:data <=32'h00790125;14'd15428:data <=32'h009500C3;
14'd15429:data <=32'h00A200A7;14'd15430:data <=32'h00AD008F;14'd15431:data <=32'h00B2007C;
14'd15432:data <=32'h00BC0069;14'd15433:data <=32'h00C80055;14'd15434:data <=32'h00D5003E;
14'd15435:data <=32'h00DE001F;14'd15436:data <=32'h00E0FFFD;14'd15437:data <=32'h00DAFFDB;
14'd15438:data <=32'h00CCFFBB;14'd15439:data <=32'h00BAFFA0;14'd15440:data <=32'h00A3FF8A;
14'd15441:data <=32'h008AFF78;14'd15442:data <=32'h0070FF6C;14'd15443:data <=32'h0053FF63;
14'd15444:data <=32'h0035FF5E;14'd15445:data <=32'h0014FF63;14'd15446:data <=32'hFFF7FF6F;
14'd15447:data <=32'hFFDDFF84;14'd15448:data <=32'hFFCBFFA0;14'd15449:data <=32'hFFC6FFC0;
14'd15450:data <=32'hFFCCFFDD;14'd15451:data <=32'hFFDDFFF4;14'd15452:data <=32'hFFF40001;
14'd15453:data <=32'h000C0002;14'd15454:data <=32'h0021FFF9;14'd15455:data <=32'h002FFFE9;
14'd15456:data <=32'h0035FFD5;14'd15457:data <=32'h0034FFC2;14'd15458:data <=32'h002CFFB2;
14'd15459:data <=32'h0020FFA5;14'd15460:data <=32'h0013FF9D;14'd15461:data <=32'h0003FF98;
14'd15462:data <=32'hFFF5FF96;14'd15463:data <=32'hFFE5FF97;14'd15464:data <=32'hFFD8FF9D;
14'd15465:data <=32'hFFCBFFA6;14'd15466:data <=32'hFFC3FFB1;14'd15467:data <=32'hFFC1FFBE;
14'd15468:data <=32'hFFC4FFC9;14'd15469:data <=32'hFFCAFFCD;14'd15470:data <=32'hFFD1FFCE;
14'd15471:data <=32'hFFD7FFC5;14'd15472:data <=32'hFFD6FFB7;14'd15473:data <=32'hFFCCFFA9;
14'd15474:data <=32'hFFB9FF9C;14'd15475:data <=32'hFF9FFF98;14'd15476:data <=32'hFF80FF9C;
14'd15477:data <=32'hFF64FFAB;14'd15478:data <=32'hFF4DFFC4;14'd15479:data <=32'hFF3DFFE2;
14'd15480:data <=32'hFF340001;14'd15481:data <=32'hFF330021;14'd15482:data <=32'hFF360040;
14'd15483:data <=32'hFF3E005C;14'd15484:data <=32'hFF4A0079;14'd15485:data <=32'hFF590092;
14'd15486:data <=32'hFF6F00AB;14'd15487:data <=32'hFF8A00BF;14'd15488:data <=32'hFF340108;
14'd15489:data <=32'hFF650141;14'd15490:data <=32'hFF9A0150;14'd15491:data <=32'hFF9800C4;
14'd15492:data <=32'hFFA2008B;14'd15493:data <=32'hFFA5009B;14'd15494:data <=32'hFFAD00B3;
14'd15495:data <=32'hFFBA00CF;14'd15496:data <=32'hFFD600EB;14'd15497:data <=32'hFFFE0103;
14'd15498:data <=32'h0030010E;14'd15499:data <=32'h0066010B;14'd15500:data <=32'h009C00F7;
14'd15501:data <=32'h00CB00D6;14'd15502:data <=32'h00EF00AA;14'd15503:data <=32'h01070078;
14'd15504:data <=32'h01120043;14'd15505:data <=32'h0114000D;14'd15506:data <=32'h0109FFDA;
14'd15507:data <=32'h00F2FFAB;14'd15508:data <=32'h00D2FF81;14'd15509:data <=32'h00A7FF62;
14'd15510:data <=32'h0075FF4F;14'd15511:data <=32'h0043FF4C;14'd15512:data <=32'h0013FF59;
14'd15513:data <=32'hFFEDFF73;14'd15514:data <=32'hFFD3FF96;14'd15515:data <=32'hFFC8FFBC;
14'd15516:data <=32'hFFCBFFDF;14'd15517:data <=32'hFFD9FFFA;14'd15518:data <=32'hFFED000D;
14'd15519:data <=32'h00020017;14'd15520:data <=32'h00160018;14'd15521:data <=32'h00270016;
14'd15522:data <=32'h0036000F;14'd15523:data <=32'h00440008;14'd15524:data <=32'h004FFFFC;
14'd15525:data <=32'h0059FFEE;14'd15526:data <=32'h0060FFDD;14'd15527:data <=32'h0063FFCA;
14'd15528:data <=32'h0061FFB4;14'd15529:data <=32'h0059FFA1;14'd15530:data <=32'h004FFF8F;
14'd15531:data <=32'h0040FF80;14'd15532:data <=32'h0031FF74;14'd15533:data <=32'h0020FF6B;
14'd15534:data <=32'h0011FF62;14'd15535:data <=32'hFFFFFF59;14'd15536:data <=32'hFFE8FF51;
14'd15537:data <=32'hFFCEFF4B;14'd15538:data <=32'hFFAFFF4B;14'd15539:data <=32'hFF8DFF53;
14'd15540:data <=32'hFF6CFF65;14'd15541:data <=32'hFF50FF82;14'd15542:data <=32'hFF3DFFA4;
14'd15543:data <=32'hFF36FFCB;14'd15544:data <=32'hFF3AFFF0;14'd15545:data <=32'hFF47000E;
14'd15546:data <=32'hFF5A0025;14'd15547:data <=32'hFF6D0033;14'd15548:data <=32'hFF7E003A;
14'd15549:data <=32'hFF8D003D;14'd15550:data <=32'hFF99003D;14'd15551:data <=32'hFFA10039;
14'd15552:data <=32'hFEE9001B;14'd15553:data <=32'hFEDF0059;14'd15554:data <=32'hFF01008C;
14'd15555:data <=32'hFF9B004C;14'd15556:data <=32'hFF940004;14'd15557:data <=32'hFF7B000A;
14'd15558:data <=32'hFF62001E;14'd15559:data <=32'hFF4E003D;14'd15560:data <=32'hFF460068;
14'd15561:data <=32'hFF4E0097;14'd15562:data <=32'hFF6600C5;14'd15563:data <=32'hFF8C00EA;
14'd15564:data <=32'hFFBB0103;14'd15565:data <=32'hFFEE010E;14'd15566:data <=32'h0022010A;
14'd15567:data <=32'h005100FC;14'd15568:data <=32'h007A00E6;14'd15569:data <=32'h009E00C7;
14'd15570:data <=32'h00BA00A4;14'd15571:data <=32'h00CE007B;14'd15572:data <=32'h00D9004F;
14'd15573:data <=32'h00D80021;14'd15574:data <=32'h00CAFFF8;14'd15575:data <=32'h00B3FFD4;
14'd15576:data <=32'h0095FFBA;14'd15577:data <=32'h0073FFAD;14'd15578:data <=32'h0054FFAB;
14'd15579:data <=32'h003AFFB0;14'd15580:data <=32'h0028FFBA;14'd15581:data <=32'h001AFFC5;
14'd15582:data <=32'h0012FFCF;14'd15583:data <=32'h000AFFD8;14'd15584:data <=32'h0003FFE2;
14'd15585:data <=32'hFFFCFFEC;14'd15586:data <=32'hFFF8FFFB;14'd15587:data <=32'hFFF9000D;
14'd15588:data <=32'hFFFE0020;14'd15589:data <=32'h000D0031;14'd15590:data <=32'h0023003F;
14'd15591:data <=32'h003D0045;14'd15592:data <=32'h005A0042;14'd15593:data <=32'h00760036;
14'd15594:data <=32'h00900022;14'd15595:data <=32'h00A40009;14'd15596:data <=32'h00B5FFE9;
14'd15597:data <=32'h00BDFFC5;14'd15598:data <=32'h00BEFF9E;14'd15599:data <=32'h00B7FF73;
14'd15600:data <=32'h00A5FF47;14'd15601:data <=32'h0085FF1E;14'd15602:data <=32'h005AFEFD;
14'd15603:data <=32'h0025FEE6;14'd15604:data <=32'hFFEBFEE1;14'd15605:data <=32'hFFAEFEEC;
14'd15606:data <=32'hFF79FF07;14'd15607:data <=32'hFF50FF30;14'd15608:data <=32'hFF36FF5E;
14'd15609:data <=32'hFF2CFF8E;14'd15610:data <=32'hFF2EFFB9;14'd15611:data <=32'hFF3AFFDE;
14'd15612:data <=32'hFF4AFFF9;14'd15613:data <=32'hFF5E000C;14'd15614:data <=32'hFF710019;
14'd15615:data <=32'hFF83001F;14'd15616:data <=32'hFF74FFBE;14'd15617:data <=32'hFF5EFFC7;
14'd15618:data <=32'hFF4EFFED;14'd15619:data <=32'hFF6A003B;14'd15620:data <=32'hFF77FFF8;
14'd15621:data <=32'hFF6FFFFC;14'd15622:data <=32'hFF650007;14'd15623:data <=32'hFF590016;
14'd15624:data <=32'hFF500030;14'd15625:data <=32'hFF51004E;14'd15626:data <=32'hFF5C006E;
14'd15627:data <=32'hFF710089;14'd15628:data <=32'hFF8D009E;14'd15629:data <=32'hFFAA00A8;
14'd15630:data <=32'hFFC800AA;14'd15631:data <=32'hFFE000A7;14'd15632:data <=32'hFFF4009F;
14'd15633:data <=32'h00050099;14'd15634:data <=32'h00140091;14'd15635:data <=32'h0023008A;
14'd15636:data <=32'h002F0080;14'd15637:data <=32'h003B0074;14'd15638:data <=32'h00440066;
14'd15639:data <=32'h0048005A;14'd15640:data <=32'h0049004F;14'd15641:data <=32'h004A0047;
14'd15642:data <=32'h004A0041;14'd15643:data <=32'h004F003D;14'd15644:data <=32'h00550036;
14'd15645:data <=32'h005D002C;14'd15646:data <=32'h0062001D;14'd15647:data <=32'h0062000A;
14'd15648:data <=32'h005BFFF6;14'd15649:data <=32'h004BFFE4;14'd15650:data <=32'h0036FFDB;
14'd15651:data <=32'h001DFFDB;14'd15652:data <=32'h0007FFE4;14'd15653:data <=32'hFFF5FFF7;
14'd15654:data <=32'hFFED000F;14'd15655:data <=32'hFFEE002A;14'd15656:data <=32'hFFFA0043;
14'd15657:data <=32'h000E0057;14'd15658:data <=32'h00280066;14'd15659:data <=32'h0046006D;
14'd15660:data <=32'h0067006C;14'd15661:data <=32'h008A0063;14'd15662:data <=32'h00AC004F;
14'd15663:data <=32'h00CB0032;14'd15664:data <=32'h00E30009;14'd15665:data <=32'h00F0FFDA;
14'd15666:data <=32'h00EFFFA7;14'd15667:data <=32'h00E0FF72;14'd15668:data <=32'h00C3FF45;
14'd15669:data <=32'h009AFF23;14'd15670:data <=32'h006DFF0D;14'd15671:data <=32'h003FFF06;
14'd15672:data <=32'h0015FF09;14'd15673:data <=32'hFFF3FF13;14'd15674:data <=32'hFFD7FF21;
14'd15675:data <=32'hFFBFFF2D;14'd15676:data <=32'hFFABFF3B;14'd15677:data <=32'hFF98FF47;
14'd15678:data <=32'hFF85FF55;14'd15679:data <=32'hFF73FF65;14'd15680:data <=32'hFF8BFFD1;
14'd15681:data <=32'hFF90FFD3;14'd15682:data <=32'hFF87FFC9;14'd15683:data <=32'hFF36FF7F;
14'd15684:data <=32'hFF2BFF58;14'd15685:data <=32'hFF12FF79;14'd15686:data <=32'hFEFDFFA0;
14'd15687:data <=32'hFEEFFFCD;14'd15688:data <=32'hFEEBFFFE;14'd15689:data <=32'hFEF30033;
14'd15690:data <=32'hFF0B0064;14'd15691:data <=32'hFF2E008D;14'd15692:data <=32'hFF5D00A8;
14'd15693:data <=32'hFF8E00B4;14'd15694:data <=32'hFFBB00AF;14'd15695:data <=32'hFFE000A0;
14'd15696:data <=32'hFFFA0088;14'd15697:data <=32'h00090070;14'd15698:data <=32'h000F0058;
14'd15699:data <=32'h000E0044;14'd15700:data <=32'h00080036;14'd15701:data <=32'h0001002C;
14'd15702:data <=32'hFFF60025;14'd15703:data <=32'hFFEA0023;14'd15704:data <=32'hFFDF0028;
14'd15705:data <=32'hFFD50032;14'd15706:data <=32'hFFD00042;14'd15707:data <=32'hFFD40055;
14'd15708:data <=32'hFFDF0066;14'd15709:data <=32'hFFF30073;14'd15710:data <=32'h000A0078;
14'd15711:data <=32'h00230073;14'd15712:data <=32'h00360064;14'd15713:data <=32'h00410050;
14'd15714:data <=32'h0045003C;14'd15715:data <=32'h00400029;14'd15716:data <=32'h0036001E;
14'd15717:data <=32'h002A0019;14'd15718:data <=32'h001D001B;14'd15719:data <=32'h00150021;
14'd15720:data <=32'h00110029;14'd15721:data <=32'h00110033;14'd15722:data <=32'h0014003C;
14'd15723:data <=32'h001A0044;14'd15724:data <=32'h0023004D;14'd15725:data <=32'h002F0055;
14'd15726:data <=32'h003E005B;14'd15727:data <=32'h0051005D;14'd15728:data <=32'h0067005A;
14'd15729:data <=32'h007D0050;14'd15730:data <=32'h00910040;14'd15731:data <=32'h00A0002B;
14'd15732:data <=32'h00A80016;14'd15733:data <=32'h00AC0000;14'd15734:data <=32'h00ACFFEC;
14'd15735:data <=32'h00ACFFDC;14'd15736:data <=32'h00ADFFCC;14'd15737:data <=32'h00B1FFBB;
14'd15738:data <=32'h00B6FFA5;14'd15739:data <=32'h00BAFF89;14'd15740:data <=32'h00B7FF64;
14'd15741:data <=32'h00AAFF3C;14'd15742:data <=32'h0091FF16;14'd15743:data <=32'h006BFEF3;
14'd15744:data <=32'hFFBAFF65;14'd15745:data <=32'hFFB6FF6D;14'd15746:data <=32'hFFC7FF69;
14'd15747:data <=32'h001AFEE6;14'd15748:data <=32'hFFEDFE9B;14'd15749:data <=32'hFFA8FEA2;
14'd15750:data <=32'hFF65FEB7;14'd15751:data <=32'hFF28FEDC;14'd15752:data <=32'hFEF5FF11;
14'd15753:data <=32'hFECFFF52;14'd15754:data <=32'hFEBEFF9C;14'd15755:data <=32'hFEC1FFE5;
14'd15756:data <=32'hFEDA0026;14'd15757:data <=32'hFF010059;14'd15758:data <=32'hFF30007C;
14'd15759:data <=32'hFF61008D;14'd15760:data <=32'hFF8E0090;14'd15761:data <=32'hFFB40089;
14'd15762:data <=32'hFFD1007C;14'd15763:data <=32'hFFE7006B;14'd15764:data <=32'hFFF70058;
14'd15765:data <=32'h00010045;14'd15766:data <=32'h00040031;14'd15767:data <=32'h0001001F;
14'd15768:data <=32'hFFF80010;14'd15769:data <=32'hFFEB0007;14'd15770:data <=32'hFFDC0005;
14'd15771:data <=32'hFFCC000A;14'd15772:data <=32'hFFC30014;14'd15773:data <=32'hFFBF0022;
14'd15774:data <=32'hFFC1002F;14'd15775:data <=32'hFFC70039;14'd15776:data <=32'hFFCD003F;
14'd15777:data <=32'hFFD50042;14'd15778:data <=32'hFFD80042;14'd15779:data <=32'hFFD80044;
14'd15780:data <=32'hFFD6004A;14'd15781:data <=32'hFFD70053;14'd15782:data <=32'hFFDB005F;
14'd15783:data <=32'hFFE4006C;14'd15784:data <=32'hFFF30076;14'd15785:data <=32'h0005007B;
14'd15786:data <=32'h00180079;14'd15787:data <=32'h002A0074;14'd15788:data <=32'h0038006A;
14'd15789:data <=32'h0042005E;14'd15790:data <=32'h00480053;14'd15791:data <=32'h004B0049;
14'd15792:data <=32'h004C003F;14'd15793:data <=32'h004C0037;14'd15794:data <=32'h004B0030;
14'd15795:data <=32'h0046002C;14'd15796:data <=32'h0041002B;14'd15797:data <=32'h003B002E;
14'd15798:data <=32'h00380038;14'd15799:data <=32'h003C0047;14'd15800:data <=32'h0049005A;
14'd15801:data <=32'h00630067;14'd15802:data <=32'h0087006D;14'd15803:data <=32'h00B10066;
14'd15804:data <=32'h00DC004E;14'd15805:data <=32'h01020026;14'd15806:data <=32'h011AFFF2;
14'd15807:data <=32'h0125FFB5;14'd15808:data <=32'h0093FF8B;14'd15809:data <=32'h0096FF6F;
14'd15810:data <=32'h009CFF6D;14'd15811:data <=32'h00E4FF86;14'd15812:data <=32'h00DAFF15;
14'd15813:data <=32'h00ADFEEF;14'd15814:data <=32'h0077FED1;14'd15815:data <=32'h003CFEC1;
14'd15816:data <=32'hFFFDFEBF;14'd15817:data <=32'hFFC1FECE;14'd15818:data <=32'hFF8CFEED;
14'd15819:data <=32'hFF64FF16;14'd15820:data <=32'hFF4BFF43;14'd15821:data <=32'hFF41FF70;
14'd15822:data <=32'hFF40FF97;14'd15823:data <=32'hFF45FFB7;14'd15824:data <=32'hFF4EFFD1;
14'd15825:data <=32'hFF56FFE7;14'd15826:data <=32'hFF5EFFF9;14'd15827:data <=32'hFF66000C;
14'd15828:data <=32'hFF72001F;14'd15829:data <=32'hFF81002E;14'd15830:data <=32'hFF94003A;
14'd15831:data <=32'hFFA70041;14'd15832:data <=32'hFFBA0042;14'd15833:data <=32'hFFCB003F;
14'd15834:data <=32'hFFD80039;14'd15835:data <=32'hFFE10032;14'd15836:data <=32'hFFE9002B;
14'd15837:data <=32'hFFF00023;14'd15838:data <=32'hFFF50018;14'd15839:data <=32'hFFF7000C;
14'd15840:data <=32'hFFF6FFFC;14'd15841:data <=32'hFFEDFFED;14'd15842:data <=32'hFFDEFFE0;
14'd15843:data <=32'hFFC7FFDB;14'd15844:data <=32'hFFACFFDD;14'd15845:data <=32'hFF92FFEC;
14'd15846:data <=32'hFF7E0004;14'd15847:data <=32'hFF720024;14'd15848:data <=32'hFF730046;
14'd15849:data <=32'hFF7E0067;14'd15850:data <=32'hFF920083;14'd15851:data <=32'hFFAD0096;
14'd15852:data <=32'hFFCA00A1;14'd15853:data <=32'hFFE600A4;14'd15854:data <=32'h000100A2;
14'd15855:data <=32'h00170099;14'd15856:data <=32'h002B008D;14'd15857:data <=32'h0039007E;
14'd15858:data <=32'h0043006E;14'd15859:data <=32'h0047005D;14'd15860:data <=32'h0044004E;
14'd15861:data <=32'h003D0042;14'd15862:data <=32'h0031003F;14'd15863:data <=32'h00270046;
14'd15864:data <=32'h00220054;14'd15865:data <=32'h00270068;14'd15866:data <=32'h0037007B;
14'd15867:data <=32'h0053008A;14'd15868:data <=32'h0077008E;14'd15869:data <=32'h009E0084;
14'd15870:data <=32'h00C2006D;14'd15871:data <=32'h00DE004D;14'd15872:data <=32'h00A70081;
14'd15873:data <=32'h00E0006D;14'd15874:data <=32'h00F8004F;14'd15875:data <=32'h00B50017;
14'd15876:data <=32'h00C5FFBD;14'd15877:data <=32'h00B7FFA5;14'd15878:data <=32'h00A7FF90;
14'd15879:data <=32'h0094FF7D;14'd15880:data <=32'h007EFF6F;14'd15881:data <=32'h0066FF66;
14'd15882:data <=32'h004EFF64;14'd15883:data <=32'h003CFF66;14'd15884:data <=32'h002FFF6A;
14'd15885:data <=32'h0026FF6C;14'd15886:data <=32'h0021FF6A;14'd15887:data <=32'h0018FF61;
14'd15888:data <=32'h000BFF56;14'd15889:data <=32'hFFF5FF4B;14'd15890:data <=32'hFFD9FF46;
14'd15891:data <=32'hFFB7FF49;14'd15892:data <=32'hFF96FF56;14'd15893:data <=32'hFF7AFF6F;
14'd15894:data <=32'hFF66FF8D;14'd15895:data <=32'hFF59FFB0;14'd15896:data <=32'hFF58FFD3;
14'd15897:data <=32'hFF5EFFF2;14'd15898:data <=32'hFF6B000F;14'd15899:data <=32'hFF7D0028;
14'd15900:data <=32'hFF94003A;14'd15901:data <=32'hFFAE0046;14'd15902:data <=32'hFFCD004B;
14'd15903:data <=32'hFFEB0045;14'd15904:data <=32'h00060035;14'd15905:data <=32'h0019001B;
14'd15906:data <=32'h0020FFFD;14'd15907:data <=32'h001BFFDC;14'd15908:data <=32'h000AFFC0;
14'd15909:data <=32'hFFEEFFAD;14'd15910:data <=32'hFFCEFFA6;14'd15911:data <=32'hFFAEFFAA;
14'd15912:data <=32'hFF92FFB9;14'd15913:data <=32'hFF7CFFCE;14'd15914:data <=32'hFF6EFFE6;
14'd15915:data <=32'hFF660000;14'd15916:data <=32'hFF640018;14'd15917:data <=32'hFF650030;
14'd15918:data <=32'hFF6A0046;14'd15919:data <=32'hFF72005A;14'd15920:data <=32'hFF7C0070;
14'd15921:data <=32'hFF8A0083;14'd15922:data <=32'hFF9B0094;14'd15923:data <=32'hFFAE00A0;
14'd15924:data <=32'hFFC100A8;14'd15925:data <=32'hFFD500AE;14'd15926:data <=32'hFFE600B3;
14'd15927:data <=32'hFFF600B8;14'd15928:data <=32'h000700BF;14'd15929:data <=32'h001D00C6;
14'd15930:data <=32'h003900CC;14'd15931:data <=32'h005A00CC;14'd15932:data <=32'h008000C1;
14'd15933:data <=32'h00A300AF;14'd15934:data <=32'h00C1008F;14'd15935:data <=32'h00D40069;
14'd15936:data <=32'hFFF700BF;14'd15937:data <=32'h002D00E2;14'd15938:data <=32'h007100DF;
14'd15939:data <=32'h00B9002D;14'd15940:data <=32'h00BEFFD3;14'd15941:data <=32'h00A3FFC0;
14'd15942:data <=32'h0087FFB6;14'd15943:data <=32'h0070FFB4;14'd15944:data <=32'h0059FFB7;
14'd15945:data <=32'h0047FFC0;14'd15946:data <=32'h003CFFCD;14'd15947:data <=32'h0039FFDD;
14'd15948:data <=32'h0040FFEB;14'd15949:data <=32'h0050FFF3;14'd15950:data <=32'h0065FFF2;
14'd15951:data <=32'h007BFFE5;14'd15952:data <=32'h008BFFCA;14'd15953:data <=32'h0090FFA9;
14'd15954:data <=32'h0087FF84;14'd15955:data <=32'h0072FF64;14'd15956:data <=32'h0053FF4B;
14'd15957:data <=32'h002DFF3D;14'd15958:data <=32'h0007FF3B;14'd15959:data <=32'hFFE3FF42;
14'd15960:data <=32'hFFC4FF51;14'd15961:data <=32'hFFAAFF65;14'd15962:data <=32'hFF95FF7E;
14'd15963:data <=32'hFF88FF99;14'd15964:data <=32'hFF7FFFB7;14'd15965:data <=32'hFF80FFD6;
14'd15966:data <=32'hFF89FFF3;14'd15967:data <=32'hFF9C000C;14'd15968:data <=32'hFFB3001B;
14'd15969:data <=32'hFFCD0021;14'd15970:data <=32'hFFE5001D;14'd15971:data <=32'hFFF90011;
14'd15972:data <=32'h00050000;14'd15973:data <=32'h000AFFED;14'd15974:data <=32'h0007FFDD;
14'd15975:data <=32'h0000FFCF;14'd15976:data <=32'hFFF9FFC6;14'd15977:data <=32'hFFF0FFBE;
14'd15978:data <=32'hFFE8FFB6;14'd15979:data <=32'hFFDEFFAE;14'd15980:data <=32'hFFD0FFA5;
14'd15981:data <=32'hFFBFFF9C;14'd15982:data <=32'hFFA6FF96;14'd15983:data <=32'hFF89FF97;
14'd15984:data <=32'hFF6AFFA1;14'd15985:data <=32'hFF4BFFB3;14'd15986:data <=32'hFF2FFFCF;
14'd15987:data <=32'hFF1AFFF2;14'd15988:data <=32'hFF0D001B;14'd15989:data <=32'hFF070046;
14'd15990:data <=32'hFF090074;14'd15991:data <=32'hFF1500A4;14'd15992:data <=32'hFF2C00D5;
14'd15993:data <=32'hFF4D0102;14'd15994:data <=32'hFF7C012A;14'd15995:data <=32'hFFB60147;
14'd15996:data <=32'hFFF90154;14'd15997:data <=32'h0040014F;14'd15998:data <=32'h00820136;
14'd15999:data <=32'h00BA010C;14'd16000:data <=32'hFFD40088;14'd16001:data <=32'hFFE700B1;
14'd16002:data <=32'h001500DB;14'd16003:data <=32'h00B900D6;14'd16004:data <=32'h00DC0069;
14'd16005:data <=32'h00D4003F;14'd16006:data <=32'h00C5001D;14'd16007:data <=32'h00B30002;
14'd16008:data <=32'h009DFFEF;14'd16009:data <=32'h0085FFE2;14'd16010:data <=32'h006DFFDF;
14'd16011:data <=32'h005BFFE3;14'd16012:data <=32'h004FFFEE;14'd16013:data <=32'h004DFFFB;
14'd16014:data <=32'h00540005;14'd16015:data <=32'h00610007;14'd16016:data <=32'h00700000;
14'd16017:data <=32'h007CFFF1;14'd16018:data <=32'h0081FFDB;14'd16019:data <=32'h007EFFC5;
14'd16020:data <=32'h0073FFB1;14'd16021:data <=32'h0063FFA2;14'd16022:data <=32'h0051FF99;
14'd16023:data <=32'h0041FF96;14'd16024:data <=32'h0033FF94;14'd16025:data <=32'h0027FF94;
14'd16026:data <=32'h001CFF95;14'd16027:data <=32'h0010FF95;14'd16028:data <=32'h0004FF98;
14'd16029:data <=32'hFFF9FF9C;14'd16030:data <=32'hFFEEFFA4;14'd16031:data <=32'hFFE7FFAC;
14'd16032:data <=32'hFFE3FFB7;14'd16033:data <=32'hFFE2FFBE;14'd16034:data <=32'hFFE3FFC3;
14'd16035:data <=32'hFFE2FFC8;14'd16036:data <=32'hFFE1FFCA;14'd16037:data <=32'hFFDEFFCE;
14'd16038:data <=32'hFFDCFFD3;14'd16039:data <=32'hFFDDFFDC;14'd16040:data <=32'hFFE0FFE7;
14'd16041:data <=32'hFFEAFFEE;14'd16042:data <=32'hFFFAFFF2;14'd16043:data <=32'h000CFFEC;
14'd16044:data <=32'h001CFFDD;14'd16045:data <=32'h0027FFC5;14'd16046:data <=32'h0028FFA6;
14'd16047:data <=32'h001DFF86;14'd16048:data <=32'h0006FF68;14'd16049:data <=32'hFFE4FF51;
14'd16050:data <=32'hFFBAFF44;14'd16051:data <=32'hFF8CFF43;14'd16052:data <=32'hFF5DFF4D;
14'd16053:data <=32'hFF30FF64;14'd16054:data <=32'hFF05FF84;14'd16055:data <=32'hFEE1FFB1;
14'd16056:data <=32'hFEC5FFE8;14'd16057:data <=32'hFEB80028;14'd16058:data <=32'hFEBB006C;
14'd16059:data <=32'hFED000B0;14'd16060:data <=32'hFEF800ED;14'd16061:data <=32'hFF30011C;
14'd16062:data <=32'hFF71013B;14'd16063:data <=32'hFFB50146;14'd16064:data <=32'hFF9F00CD;
14'd16065:data <=32'hFFB800EB;14'd16066:data <=32'hFFC6010B;14'd16067:data <=32'hFFC10131;
14'd16068:data <=32'h000000EE;14'd16069:data <=32'h001B00E6;14'd16070:data <=32'h003500DD;
14'd16071:data <=32'h004E00D2;14'd16072:data <=32'h006600C1;14'd16073:data <=32'h007A00AF;
14'd16074:data <=32'h008A0098;14'd16075:data <=32'h00960083;14'd16076:data <=32'h009F006F;
14'd16077:data <=32'h00A8005B;14'd16078:data <=32'h00B00046;14'd16079:data <=32'h00B7002E;
14'd16080:data <=32'h00BC0012;14'd16081:data <=32'h00B8FFF2;14'd16082:data <=32'h00AEFFD3;
14'd16083:data <=32'h0098FFB7;14'd16084:data <=32'h007CFFA3;14'd16085:data <=32'h005CFF9A;
14'd16086:data <=32'h003CFF9D;14'd16087:data <=32'h0022FFA9;14'd16088:data <=32'h0011FFBB;
14'd16089:data <=32'h000AFFCF;14'd16090:data <=32'h000DFFE0;14'd16091:data <=32'h0012FFED;
14'd16092:data <=32'h001CFFF5;14'd16093:data <=32'h0026FFF8;14'd16094:data <=32'h0030FFF7;
14'd16095:data <=32'h003AFFF3;14'd16096:data <=32'h0043FFEB;14'd16097:data <=32'h0049FFE1;
14'd16098:data <=32'h004DFFD3;14'd16099:data <=32'h004BFFC2;14'd16100:data <=32'h0044FFB1;
14'd16101:data <=32'h0036FFA4;14'd16102:data <=32'h0023FF9D;14'd16103:data <=32'h0012FF9D;
14'd16104:data <=32'h0000FFA6;14'd16105:data <=32'hFFF5FFB3;14'd16106:data <=32'hFFF4FFC2;
14'd16107:data <=32'hFFFAFFCF;14'd16108:data <=32'h0007FFD5;14'd16109:data <=32'h0017FFD2;
14'd16110:data <=32'h0024FFC7;14'd16111:data <=32'h002DFFB3;14'd16112:data <=32'h002BFF9D;
14'd16113:data <=32'h0021FF85;14'd16114:data <=32'h0011FF71;14'd16115:data <=32'hFFFBFF60;
14'd16116:data <=32'hFFE0FF55;14'd16117:data <=32'hFFC2FF4E;14'd16118:data <=32'hFFA2FF4E;
14'd16119:data <=32'hFF7FFF54;14'd16120:data <=32'hFF5CFF63;14'd16121:data <=32'hFF3CFF7C;
14'd16122:data <=32'hFF1FFF9C;14'd16123:data <=32'hFF0CFFC3;14'd16124:data <=32'hFF04FFF0;
14'd16125:data <=32'hFF07001A;14'd16126:data <=32'hFF14003F;14'd16127:data <=32'hFF27005D;
14'd16128:data <=32'hFEE1007E;14'd16129:data <=32'hFEEF00B6;14'd16130:data <=32'hFF0600D0;
14'd16131:data <=32'hFF1A005C;14'd16132:data <=32'hFF340039;14'd16133:data <=32'hFF2D005A;
14'd16134:data <=32'hFF2F0080;14'd16135:data <=32'hFF3B00AC;14'd16136:data <=32'hFF5400D3;
14'd16137:data <=32'hFF7800F3;14'd16138:data <=32'hFFA1010E;14'd16139:data <=32'hFFCF011C;
14'd16140:data <=32'h00010123;14'd16141:data <=32'h00350120;14'd16142:data <=32'h00690113;
14'd16143:data <=32'h009B00F8;14'd16144:data <=32'h00C600D0;14'd16145:data <=32'h00E7009F;
14'd16146:data <=32'h00F90064;14'd16147:data <=32'h00F90028;14'd16148:data <=32'h00E7FFF0;
14'd16149:data <=32'h00C7FFC3;14'd16150:data <=32'h009CFFA6;14'd16151:data <=32'h0070FF98;
14'd16152:data <=32'h0046FF98;14'd16153:data <=32'h0024FFA4;14'd16154:data <=32'h000BFFB7;
14'd16155:data <=32'hFFFBFFCD;14'd16156:data <=32'hFFF3FFE3;14'd16157:data <=32'hFFF1FFF9;
14'd16158:data <=32'hFFF5000C;14'd16159:data <=32'hFFFE001F;14'd16160:data <=32'h000D002D;
14'd16161:data <=32'h00200036;14'd16162:data <=32'h00350038;14'd16163:data <=32'h004B0034;
14'd16164:data <=32'h005D0027;14'd16165:data <=32'h006A0016;14'd16166:data <=32'h00700004;
14'd16167:data <=32'h0071FFF2;14'd16168:data <=32'h006FFFE4;14'd16169:data <=32'h006CFFD8;
14'd16170:data <=32'h0068FFCE;14'd16171:data <=32'h0069FFC7;14'd16172:data <=32'h006AFFBC;
14'd16173:data <=32'h006BFFAC;14'd16174:data <=32'h006AFF98;14'd16175:data <=32'h0062FF83;
14'd16176:data <=32'h0053FF6D;14'd16177:data <=32'h003DFF5B;14'd16178:data <=32'h0022FF4F;
14'd16179:data <=32'h0004FF4B;14'd16180:data <=32'hFFE9FF4E;14'd16181:data <=32'hFFD0FF58;
14'd16182:data <=32'hFFBCFF63;14'd16183:data <=32'hFFACFF70;14'd16184:data <=32'hFF9FFF7F;
14'd16185:data <=32'hFF94FF8F;14'd16186:data <=32'hFF8CFF9F;14'd16187:data <=32'hFF89FFB0;
14'd16188:data <=32'hFF8AFFBF;14'd16189:data <=32'hFF8FFFCB;14'd16190:data <=32'hFF96FFD1;
14'd16191:data <=32'hFF9CFFCF;14'd16192:data <=32'hFF03FF86;14'd16193:data <=32'hFEE1FFAE;
14'd16194:data <=32'hFEE5FFDB;14'd16195:data <=32'hFF7BFFC4;14'd16196:data <=32'hFF80FF86;
14'd16197:data <=32'hFF58FF8E;14'd16198:data <=32'hFF30FFA6;14'd16199:data <=32'hFF10FFCA;
14'd16200:data <=32'hFEFCFFF9;14'd16201:data <=32'hFEF4002B;14'd16202:data <=32'hFEF9005E;
14'd16203:data <=32'hFF090090;14'd16204:data <=32'hFF2400BD;14'd16205:data <=32'hFF4800E4;
14'd16206:data <=32'hFF760106;14'd16207:data <=32'hFFAD011B;14'd16208:data <=32'hFFE70122;
14'd16209:data <=32'h00230117;14'd16210:data <=32'h005900FE;14'd16211:data <=32'h008400D8;
14'd16212:data <=32'h009F00A9;14'd16213:data <=32'h00AA0079;14'd16214:data <=32'h00A9004E;
14'd16215:data <=32'h009D0029;14'd16216:data <=32'h008B000F;14'd16217:data <=32'h0077FFFB;
14'd16218:data <=32'h0064FFEE;14'd16219:data <=32'h0052FFE5;14'd16220:data <=32'h0040FFDF;
14'd16221:data <=32'h002EFFDC;14'd16222:data <=32'h001BFFDE;14'd16223:data <=32'h000AFFE5;
14'd16224:data <=32'hFFFBFFF1;14'd16225:data <=32'hFFF00002;14'd16226:data <=32'hFFEC0016;
14'd16227:data <=32'hFFEE002A;14'd16228:data <=32'hFFF6003B;14'd16229:data <=32'h00020049;
14'd16230:data <=32'h00110056;14'd16231:data <=32'h0023005F;14'd16232:data <=32'h00360067;
14'd16233:data <=32'h004E006B;14'd16234:data <=32'h0069006A;14'd16235:data <=32'h00890064;
14'd16236:data <=32'h00A90053;14'd16237:data <=32'h00C80038;14'd16238:data <=32'h00E00011;
14'd16239:data <=32'h00EDFFE3;14'd16240:data <=32'h00EDFFAF;14'd16241:data <=32'h00DDFF7D;
14'd16242:data <=32'h00C0FF50;14'd16243:data <=32'h0098FF2E;14'd16244:data <=32'h006AFF1A;
14'd16245:data <=32'h003CFF14;14'd16246:data <=32'h0010FF17;14'd16247:data <=32'hFFEAFF24;
14'd16248:data <=32'hFFCBFF36;14'd16249:data <=32'hFFB2FF4F;14'd16250:data <=32'hFFA0FF6A;
14'd16251:data <=32'hFF96FF86;14'd16252:data <=32'hFF96FFA1;14'd16253:data <=32'hFF9EFFBA;
14'd16254:data <=32'hFFAEFFCA;14'd16255:data <=32'hFFC2FFCF;14'd16256:data <=32'hFFCCFF6D;
14'd16257:data <=32'hFFB7FF5E;14'd16258:data <=32'hFF98FF6C;14'd16259:data <=32'hFF9DFFBB;
14'd16260:data <=32'hFFB4FF7A;14'd16261:data <=32'hFF99FF77;14'd16262:data <=32'hFF7DFF7E;
14'd16263:data <=32'hFF60FF8F;14'd16264:data <=32'hFF4BFFA7;14'd16265:data <=32'hFF3DFFC4;
14'd16266:data <=32'hFF35FFE3;14'd16267:data <=32'hFF330001;14'd16268:data <=32'hFF37001E;
14'd16269:data <=32'hFF3D003A;14'd16270:data <=32'hFF490055;14'd16271:data <=32'hFF5B006F;
14'd16272:data <=32'hFF730085;14'd16273:data <=32'hFF8E0094;14'd16274:data <=32'hFFAD009B;
14'd16275:data <=32'hFFC9009A;14'd16276:data <=32'hFFDF0092;14'd16277:data <=32'hFFEF0087;
14'd16278:data <=32'hFFFA007D;14'd16279:data <=32'h00010077;14'd16280:data <=32'h00070074;
14'd16281:data <=32'h00110074;14'd16282:data <=32'h001E0072;14'd16283:data <=32'h002D006B;
14'd16284:data <=32'h003D005F;14'd16285:data <=32'h0049004E;14'd16286:data <=32'h004E0037;
14'd16287:data <=32'h004D0022;14'd16288:data <=32'h0043000D;14'd16289:data <=32'h0035FFFE;
14'd16290:data <=32'h0022FFF6;14'd16291:data <=32'h000EFFF4;14'd16292:data <=32'hFFFBFFF8;
14'd16293:data <=32'hFFEA0003;14'd16294:data <=32'hFFDC0013;14'd16295:data <=32'hFFD10027;
14'd16296:data <=32'hFFCB0042;14'd16297:data <=32'hFFCF0060;14'd16298:data <=32'hFFDC007F;
14'd16299:data <=32'hFFF6009C;14'd16300:data <=32'h001C00B2;14'd16301:data <=32'h004900BD;
14'd16302:data <=32'h007A00B8;14'd16303:data <=32'h00AB00A5;14'd16304:data <=32'h00D40082;
14'd16305:data <=32'h00F10055;14'd16306:data <=32'h01010024;14'd16307:data <=32'h0101FFF2;
14'd16308:data <=32'h00F7FFC5;14'd16309:data <=32'h00E4FF9E;14'd16310:data <=32'h00CEFF7F;
14'd16311:data <=32'h00B3FF66;14'd16312:data <=32'h0097FF53;14'd16313:data <=32'h007AFF44;
14'd16314:data <=32'h005BFF3B;14'd16315:data <=32'h003EFF3A;14'd16316:data <=32'h0023FF3D;
14'd16317:data <=32'h000CFF46;14'd16318:data <=32'hFFFCFF4F;14'd16319:data <=32'hFFF1FF59;
14'd16320:data <=32'hFFE8FFBF;14'd16321:data <=32'hFFFDFFB6;14'd16322:data <=32'hFFFDFF9B;
14'd16323:data <=32'hFFC1FF37;14'd16324:data <=32'hFFC3FF02;14'd16325:data <=32'hFF96FF0D;
14'd16326:data <=32'hFF6CFF26;14'd16327:data <=32'hFF47FF48;14'd16328:data <=32'hFF2FFF73;
14'd16329:data <=32'hFF27FFA2;14'd16330:data <=32'hFF29FFCE;14'd16331:data <=32'hFF36FFF3;
14'd16332:data <=32'hFF490010;14'd16333:data <=32'hFF5F0026;14'd16334:data <=32'hFF760035;
14'd16335:data <=32'hFF8C003E;14'd16336:data <=32'hFFA10041;14'd16337:data <=32'hFFB6003F;
14'd16338:data <=32'hFFC80037;14'd16339:data <=32'hFFD3002A;14'd16340:data <=32'hFFD5001A;
14'd16341:data <=32'hFFD0000D;14'd16342:data <=32'hFFC30005;14'd16343:data <=32'hFFB30006;
14'd16344:data <=32'hFFA20010;14'd16345:data <=32'hFF980024;14'd16346:data <=32'hFF96003C;
14'd16347:data <=32'hFF9F0054;14'd16348:data <=32'hFFB10067;14'd16349:data <=32'hFFC80072;
14'd16350:data <=32'hFFE00075;14'd16351:data <=32'hFFF60070;14'd16352:data <=32'h00080064;
14'd16353:data <=32'h00140056;14'd16354:data <=32'h00190047;14'd16355:data <=32'h001B0038;
14'd16356:data <=32'h0019002B;14'd16357:data <=32'h00120020;14'd16358:data <=32'h00070017;
14'd16359:data <=32'hFFFB0013;14'd16360:data <=32'hFFEA0015;14'd16361:data <=32'hFFDA001F;
14'd16362:data <=32'hFFCD002F;14'd16363:data <=32'hFFC70046;14'd16364:data <=32'hFFCA005F;
14'd16365:data <=32'hFFD70079;14'd16366:data <=32'hFFEC008E;14'd16367:data <=32'h0006009A;
14'd16368:data <=32'h0022009F;14'd16369:data <=32'h003F009D;14'd16370:data <=32'h00560093;
14'd16371:data <=32'h0069008A;14'd16372:data <=32'h0079007F;14'd16373:data <=32'h00890076;
14'd16374:data <=32'h009B006B;14'd16375:data <=32'h00AE0060;14'd16376:data <=32'h00C30050;
14'd16377:data <=32'h00D70038;14'd16378:data <=32'h00EA001B;14'd16379:data <=32'h00F5FFF8;
14'd16380:data <=32'h00FBFFD3;14'd16381:data <=32'h00FBFFAD;14'd16382:data <=32'h00F2FF85;
14'd16383:data <=32'h00E6FF5E;
        
        endcase
        
end    
    
    assign dout = data;
    
endmodule
