`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 05/23/2023 02:45:31 PM
// Design Name: 
// Module Name: rom
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module sp_rom #(
    parameter integer ADDRW = 14,
    parameter integer DATA_WIDTH = 32,
    parameter RAM_TYPE = "block"
)
(
input [ADDRW-1:0] addr,
input clk,
input en,
output wire [DATA_WIDTH-1:0] dout
    );
    
//DD clock
//(*ram_style = "registers"*)reg r_clk50=0;

//wire w_xor_clk50=(r_clk50 ^ clk);

//always@(posedge w_xor_clk50) begin

//    r_clk50=~r_clk50;

//    // your code on both neg/pos
//end
 
    
 (*rom_style = RAM_TYPE*) reg [DATA_WIDTH-1:0] data;   
    
always@(negedge clk)
begin
    if(en)
    case (addr)
14'd0:data <=32'h00000000;14'd1:data <=32'h006BFFDE;14'd2:data <=32'h00BCFFB2;
14'd3:data <=32'h00D5FFA6;14'd4:data <=32'h00B8FFA4;14'd5:data <=32'h00AFFF89;
14'd6:data <=32'h00A4FF6D;14'd7:data <=32'h0095FF57;14'd8:data <=32'h0080FF39;
14'd9:data <=32'h005FFF1D;14'd10:data <=32'h0035FF0A;14'd11:data <=32'h0006FF02;
14'd12:data <=32'hFFD3FF07;14'd13:data <=32'hFFA5FF1B;14'd14:data <=32'hFF7FFF38;
14'd15:data <=32'hFF64FF5C;14'd16:data <=32'hFF51FF83;14'd17:data <=32'hFF4AFFAB;
14'd18:data <=32'hFF4AFFD2;14'd19:data <=32'hFF52FFF6;14'd20:data <=32'hFF620017;
14'd21:data <=32'hFF7B0032;14'd22:data <=32'hFF990044;14'd23:data <=32'hFFBA004C;
14'd24:data <=32'hFFDB0049;14'd25:data <=32'hFFF6003B;14'd26:data <=32'h00090024;
14'd27:data <=32'h0011000A;14'd28:data <=32'h000CFFF1;14'd29:data <=32'h0000FFDF;
14'd30:data <=32'hFFEDFFD4;14'd31:data <=32'hFFDBFFD1;14'd32:data <=32'hFFC9FFD6;
14'd33:data <=32'hFFBEFFDF;14'd34:data <=32'hFFB5FFEA;14'd35:data <=32'hFFB1FFF5;
14'd36:data <=32'hFFAEFFFE;14'd37:data <=32'hFFAD0007;14'd38:data <=32'hFFAD0010;
14'd39:data <=32'hFFAE001A;14'd40:data <=32'hFFB10022;14'd41:data <=32'hFFB50029;
14'd42:data <=32'hFFB80030;14'd43:data <=32'hFFBD0034;14'd44:data <=32'hFFC00037;
14'd45:data <=32'hFFC0003A;14'd46:data <=32'hFFBF003F;14'd47:data <=32'hFFBC0047;
14'd48:data <=32'hFFBB0053;14'd49:data <=32'hFFBE0063;14'd50:data <=32'hFFC80075;
14'd51:data <=32'hFFD70084;14'd52:data <=32'hFFEC008E;14'd53:data <=32'h00050091;
14'd54:data <=32'h001A008F;14'd55:data <=32'h002D0086;14'd56:data <=32'h0039007B;
14'd57:data <=32'h00420071;14'd58:data <=32'h0047006B;14'd59:data <=32'h004C0065;
14'd60:data <=32'h00530065;14'd61:data <=32'h005C0063;14'd62:data <=32'h00690060;
14'd63:data <=32'h0078005C;14'd64:data <=32'h00FB004C;14'd65:data <=32'h010F001F;
14'd66:data <=32'h0102FFF9;14'd67:data <=32'h00970049;14'd68:data <=32'h009D007A;
14'd69:data <=32'h00BF0068;14'd70:data <=32'h00E0004C;14'd71:data <=32'h00FC0025;
14'd72:data <=32'h010FFFF1;14'd73:data <=32'h0110FFB7;14'd74:data <=32'h0101FF7C;
14'd75:data <=32'h00E2FF47;14'd76:data <=32'h00B4FF1F;14'd77:data <=32'h007FFF04;
14'd78:data <=32'h0047FEF9;14'd79:data <=32'h0012FEFB;14'd80:data <=32'hFFE2FF0A;
14'd81:data <=32'hFFB7FF20;14'd82:data <=32'hFF95FF3E;14'd83:data <=32'hFF7AFF61;
14'd84:data <=32'hFF69FF88;14'd85:data <=32'hFF63FFB2;14'd86:data <=32'hFF68FFDA;
14'd87:data <=32'hFF77FFFD;14'd88:data <=32'hFF900017;14'd89:data <=32'hFFAD0026;
14'd90:data <=32'hFFCA002B;14'd91:data <=32'hFFE30026;14'd92:data <=32'hFFF5001B;
14'd93:data <=32'h0001000E;14'd94:data <=32'h00050000;14'd95:data <=32'h0008FFF4;
14'd96:data <=32'h0007FFEA;14'd97:data <=32'h0007FFE2;14'd98:data <=32'h0006FFD9;
14'd99:data <=32'h0002FFCC;14'd100:data <=32'hFFFBFFC1;14'd101:data <=32'hFFF0FFB5;
14'd102:data <=32'hFFE0FFAA;14'd103:data <=32'hFFCCFFA6;14'd104:data <=32'hFFB5FFA6;
14'd105:data <=32'hFF9EFFAE;14'd106:data <=32'hFF89FFBB;14'd107:data <=32'hFF77FFCD;
14'd108:data <=32'hFF69FFE1;14'd109:data <=32'hFF60FFF9;14'd110:data <=32'hFF590013;
14'd111:data <=32'hFF580030;14'd112:data <=32'hFF5D004E;14'd113:data <=32'hFF69006D;
14'd114:data <=32'hFF7D0088;14'd115:data <=32'hFF99009F;14'd116:data <=32'hFFBB00AD;
14'd117:data <=32'hFFDF00B0;14'd118:data <=32'h000200A7;14'd119:data <=32'h001D0094;
14'd120:data <=32'h002E007D;14'd121:data <=32'h00330064;14'd122:data <=32'h00300051;
14'd123:data <=32'h00250044;14'd124:data <=32'h0019003F;14'd125:data <=32'h000E0042;
14'd126:data <=32'h0008004B;14'd127:data <=32'h00060057;14'd128:data <=32'h003D00AA;
14'd129:data <=32'h005C00AB;14'd130:data <=32'h00700093;14'd131:data <=32'h00320054;
14'd132:data <=32'h002A0097;14'd133:data <=32'h004700A0;14'd134:data <=32'h006900A1;
14'd135:data <=32'h008E0097;14'd136:data <=32'h00B20080;14'd137:data <=32'h00CF005D;
14'd138:data <=32'h00E10033;14'd139:data <=32'h00E50006;14'd140:data <=32'h00DDFFDB;
14'd141:data <=32'h00CCFFB7;14'd142:data <=32'h00B5FF9A;14'd143:data <=32'h009BFF84;
14'd144:data <=32'h0081FF76;14'd145:data <=32'h0066FF6B;14'd146:data <=32'h004CFF65;
14'd147:data <=32'h0033FF63;14'd148:data <=32'h0018FF64;14'd149:data <=32'h0000FF6D;
14'd150:data <=32'hFFEAFF79;14'd151:data <=32'hFFDAFF8A;14'd152:data <=32'hFFD1FF9C;
14'd153:data <=32'hFFCCFFAD;14'd154:data <=32'hFFC9FFBA;14'd155:data <=32'hFFCAFFC6;
14'd156:data <=32'hFFC9FFCF;14'd157:data <=32'hFFCAFFDA;14'd158:data <=32'hFFC9FFE7;
14'd159:data <=32'hFFCDFFF3;14'd160:data <=32'hFFD60001;14'd161:data <=32'hFFE4000D;
14'd162:data <=32'hFFF80013;14'd163:data <=32'h000E0011;14'd164:data <=32'h00240005;
14'd165:data <=32'h0034FFF0;14'd166:data <=32'h003CFFD5;14'd167:data <=32'h003BFFB8;
14'd168:data <=32'h0030FF9C;14'd169:data <=32'h001CFF84;14'd170:data <=32'h0001FF71;
14'd171:data <=32'hFFE2FF67;14'd172:data <=32'hFFBFFF63;14'd173:data <=32'hFF9CFF68;
14'd174:data <=32'hFF7AFF75;14'd175:data <=32'hFF59FF8C;14'd176:data <=32'hFF3FFFAA;
14'd177:data <=32'hFF2AFFD1;14'd178:data <=32'hFF22FFFC;14'd179:data <=32'hFF250029;
14'd180:data <=32'hFF350052;14'd181:data <=32'hFF500074;14'd182:data <=32'hFF70008A;
14'd183:data <=32'hFF920094;14'd184:data <=32'hFFB10093;14'd185:data <=32'hFFC9008C;
14'd186:data <=32'hFFD80082;14'd187:data <=32'hFFE1007A;14'd188:data <=32'hFFE60075;
14'd189:data <=32'hFFE90073;14'd190:data <=32'hFFED0074;14'd191:data <=32'hFFF20077;
14'd192:data <=32'hFFE0003F;14'd193:data <=32'hFFD60051;14'd194:data <=32'hFFE10064;
14'd195:data <=32'h002A0081;14'd196:data <=32'h002200B4;14'd197:data <=32'h003A00AF;
14'd198:data <=32'h005400A6;14'd199:data <=32'h006D0099;14'd200:data <=32'h00830084;
14'd201:data <=32'h00950068;14'd202:data <=32'h009F0049;14'd203:data <=32'h009D0029;
14'd204:data <=32'h0093000E;14'd205:data <=32'h0082FFFA;14'd206:data <=32'h0070FFEF;
14'd207:data <=32'h0060FFED;14'd208:data <=32'h0056FFEF;14'd209:data <=32'h0052FFF2;
14'd210:data <=32'h0052FFF4;14'd211:data <=32'h0055FFF3;14'd212:data <=32'h0058FFEE;
14'd213:data <=32'h005BFFE6;14'd214:data <=32'h005AFFDD;14'd215:data <=32'h0059FFD4;
14'd216:data <=32'h0058FFC9;14'd217:data <=32'h0054FFBE;14'd218:data <=32'h004DFFB1;
14'd219:data <=32'h0041FFA4;14'd220:data <=32'h0030FF98;14'd221:data <=32'h001CFF92;
14'd222:data <=32'h0004FF93;14'd223:data <=32'hFFEDFF9D;14'd224:data <=32'hFFDBFFAE;
14'd225:data <=32'hFFD0FFC6;14'd226:data <=32'hFFD1FFE0;14'd227:data <=32'hFFDBFFF6;
14'd228:data <=32'hFFED0005;14'd229:data <=32'h0003000C;14'd230:data <=32'h001A0009;
14'd231:data <=32'h002DFFFF;14'd232:data <=32'h003BFFED;14'd233:data <=32'h0043FFD9;
14'd234:data <=32'h0045FFC3;14'd235:data <=32'h0041FFAC;14'd236:data <=32'h0038FF97;
14'd237:data <=32'h0029FF83;14'd238:data <=32'h0015FF71;14'd239:data <=32'hFFFCFF65;
14'd240:data <=32'hFFDEFF5D;14'd241:data <=32'hFFBFFF5E;14'd242:data <=32'hFFA0FF67;
14'd243:data <=32'hFF85FF77;14'd244:data <=32'hFF70FF8C;14'd245:data <=32'hFF62FFA4;
14'd246:data <=32'hFF5AFFBB;14'd247:data <=32'hFF54FFCE;14'd248:data <=32'hFF50FFE0;
14'd249:data <=32'hFF4BFFEF;14'd250:data <=32'hFF430003;14'd251:data <=32'hFF3C0019;
14'd252:data <=32'hFF360035;14'd253:data <=32'hFF370056;14'd254:data <=32'hFF400079;
14'd255:data <=32'hFF52009B;14'd256:data <=32'hFFEF002D;14'd257:data <=32'hFFDD0028;
14'd258:data <=32'hFFC10037;14'd259:data <=32'hFF8E00C2;14'd260:data <=32'hFF9E010A;
14'd261:data <=32'hFFD20113;14'd262:data <=32'h00060110;14'd263:data <=32'h00380102;
14'd264:data <=32'h006700E8;14'd265:data <=32'h008C00C3;14'd266:data <=32'h00A50095;
14'd267:data <=32'h00AE0064;14'd268:data <=32'h00A70036;14'd269:data <=32'h00950010;
14'd270:data <=32'h0079FFF7;14'd271:data <=32'h005CFFEB;14'd272:data <=32'h0041FFEB;
14'd273:data <=32'h002DFFF3;14'd274:data <=32'h0022FFFF;14'd275:data <=32'h001D000C;
14'd276:data <=32'h001E0018;14'd277:data <=32'h00230020;14'd278:data <=32'h002B0027;
14'd279:data <=32'h0035002B;14'd280:data <=32'h0041002A;14'd281:data <=32'h004F0026;
14'd282:data <=32'h005C001C;14'd283:data <=32'h0067000D;14'd284:data <=32'h006CFFFA;
14'd285:data <=32'h0069FFE5;14'd286:data <=32'h0061FFD2;14'd287:data <=32'h0051FFC5;
14'd288:data <=32'h0041FFBE;14'd289:data <=32'h002FFFBF;14'd290:data <=32'h0022FFC4;
14'd291:data <=32'h001BFFCD;14'd292:data <=32'h0019FFD6;14'd293:data <=32'h001BFFDC;
14'd294:data <=32'h001EFFDD;14'd295:data <=32'h0022FFDC;14'd296:data <=32'h0023FFDA;
14'd297:data <=32'h0023FFD7;14'd298:data <=32'h0022FFD5;14'd299:data <=32'h0022FFD3;
14'd300:data <=32'h0022FFD3;14'd301:data <=32'h0025FFD2;14'd302:data <=32'h0029FFCE;
14'd303:data <=32'h002DFFC7;14'd304:data <=32'h002FFFBE;14'd305:data <=32'h0030FFB1;
14'd306:data <=32'h002EFFA6;14'd307:data <=32'h0028FF99;14'd308:data <=32'h0022FF8C;
14'd309:data <=32'h001AFF7D;14'd310:data <=32'h000FFF6E;14'd311:data <=32'hFFFFFF5C;
14'd312:data <=32'hFFE8FF4A;14'd313:data <=32'hFFC7FF3A;14'd314:data <=32'hFF9EFF32;
14'd315:data <=32'hFF6EFF35;14'd316:data <=32'hFF3CFF47;14'd317:data <=32'hFF0CFF69;
14'd318:data <=32'hFEE7FF98;14'd319:data <=32'hFECEFFD1;14'd320:data <=32'hFF8F0010;
14'd321:data <=32'hFF810014;14'd322:data <=32'hFF67000E;14'd323:data <=32'hFEF00012;
14'd324:data <=32'hFEE2007B;14'd325:data <=32'hFF0300AC;14'd326:data <=32'hFF2E00D6;
14'd327:data <=32'hFF6000F1;14'd328:data <=32'hFF960102;14'd329:data <=32'hFFCF0103;
14'd330:data <=32'h000400F6;14'd331:data <=32'h002F00DB;14'd332:data <=32'h004D00B8;
14'd333:data <=32'h005D0094;14'd334:data <=32'h00610073;14'd335:data <=32'h005D0058;
14'd336:data <=32'h00560045;14'd337:data <=32'h004E0039;14'd338:data <=32'h00470030;
14'd339:data <=32'h0042002A;14'd340:data <=32'h003F0023;14'd341:data <=32'h003B001C;
14'd342:data <=32'h00350018;14'd343:data <=32'h002F0015;14'd344:data <=32'h00290015;
14'd345:data <=32'h00250017;14'd346:data <=32'h0025001A;14'd347:data <=32'h0027001D;
14'd348:data <=32'h0029001D;14'd349:data <=32'h002C001C;14'd350:data <=32'h002C001B;
14'd351:data <=32'h002D0019;14'd352:data <=32'h002D001B;14'd353:data <=32'h002E001E;
14'd354:data <=32'h00330022;14'd355:data <=32'h003C0025;14'd356:data <=32'h004A0025;
14'd357:data <=32'h0058001E;14'd358:data <=32'h00640012;14'd359:data <=32'h006CFFFE;
14'd360:data <=32'h006DFFEA;14'd361:data <=32'h0067FFD7;14'd362:data <=32'h005AFFC7;
14'd363:data <=32'h004AFFBD;14'd364:data <=32'h003AFFBA;14'd365:data <=32'h002BFFBD;
14'd366:data <=32'h0021FFC4;14'd367:data <=32'h001CFFCC;14'd368:data <=32'h001CFFD4;
14'd369:data <=32'h0020FFDC;14'd370:data <=32'h0026FFE0;14'd371:data <=32'h0030FFE2;
14'd372:data <=32'h003DFFE0;14'd373:data <=32'h004CFFD8;14'd374:data <=32'h005BFFC8;
14'd375:data <=32'h0067FFB0;14'd376:data <=32'h006CFF90;14'd377:data <=32'h0066FF6A;
14'd378:data <=32'h0051FF43;14'd379:data <=32'h002FFF20;14'd380:data <=32'h0000FF08;
14'd381:data <=32'hFFCAFEFE;14'd382:data <=32'hFF90FF05;14'd383:data <=32'hFF5CFF1A;
14'd384:data <=32'hFF98FF53;14'd385:data <=32'hFF6AFF51;14'd386:data <=32'hFF51FF54;
14'd387:data <=32'hFF61FF50;14'd388:data <=32'hFF2BFFA1;14'd389:data <=32'hFF23FFC4;
14'd390:data <=32'hFF20FFE9;14'd391:data <=32'hFF23000A;14'd392:data <=32'hFF2D002C;
14'd393:data <=32'hFF400048;14'd394:data <=32'hFF54005E;14'd395:data <=32'hFF6C006C;
14'd396:data <=32'hFF7F0075;14'd397:data <=32'hFF91007B;14'd398:data <=32'hFF9D0081;
14'd399:data <=32'hFFAA0089;14'd400:data <=32'hFFB90093;14'd401:data <=32'hFFCD009D;
14'd402:data <=32'hFFE500A5;14'd403:data <=32'h000200A6;14'd404:data <=32'h001E009E;
14'd405:data <=32'h0039008F;14'd406:data <=32'h004E0079;14'd407:data <=32'h0059005F;
14'd408:data <=32'h005F0045;14'd409:data <=32'h005C002C;14'd410:data <=32'h00540017;
14'd411:data <=32'h00490007;14'd412:data <=32'h003AFFF9;14'd413:data <=32'h0029FFF2;
14'd414:data <=32'h0015FFEE;14'd415:data <=32'h0001FFF2;14'd416:data <=32'hFFF0FFFD;
14'd417:data <=32'hFFE2000E;14'd418:data <=32'hFFDD0026;14'd419:data <=32'hFFE0003F;
14'd420:data <=32'hFFEE0056;14'd421:data <=32'h00040066;14'd422:data <=32'h0020006E;
14'd423:data <=32'h003C006C;14'd424:data <=32'h00540061;14'd425:data <=32'h0067004E;
14'd426:data <=32'h0072003A;14'd427:data <=32'h00770025;14'd428:data <=32'h00760013;
14'd429:data <=32'h00730004;14'd430:data <=32'h006EFFF9;14'd431:data <=32'h0069FFF0;
14'd432:data <=32'h0065FFEA;14'd433:data <=32'h0061FFE3;14'd434:data <=32'h005FFFDE;
14'd435:data <=32'h005CFFDB;14'd436:data <=32'h005CFFD7;14'd437:data <=32'h005EFFD3;
14'd438:data <=32'h0062FFCD;14'd439:data <=32'h0068FFC2;14'd440:data <=32'h006EFFB3;
14'd441:data <=32'h0071FF9D;14'd442:data <=32'h006BFF83;14'd443:data <=32'h005CFF68;
14'd444:data <=32'h0044FF51;14'd445:data <=32'h0026FF42;14'd446:data <=32'h0003FF3C;
14'd447:data <=32'hFFE1FF40;14'd448:data <=32'h006AFF26;14'd449:data <=32'h003EFEF6;
14'd450:data <=32'h000BFEE9;14'd451:data <=32'hFFE0FF66;14'd452:data <=32'hFFB9FF9E;
14'd453:data <=32'hFFBAFFA5;14'd454:data <=32'hFFBAFFA9;14'd455:data <=32'hFFB7FFA9;
14'd456:data <=32'hFFB0FFAA;14'd457:data <=32'hFFAAFFAB;14'd458:data <=32'hFFA1FFAC;
14'd459:data <=32'hFF96FFAD;14'd460:data <=32'hFF87FFAF;14'd461:data <=32'hFF73FFB6;
14'd462:data <=32'hFF5CFFC4;14'd463:data <=32'hFF47FFDC;14'd464:data <=32'hFF37FFFD;
14'd465:data <=32'hFF300026;14'd466:data <=32'hFF390052;14'd467:data <=32'hFF4D007A;
14'd468:data <=32'hFF6D009B;14'd469:data <=32'hFF9400B0;14'd470:data <=32'hFFBF00B9;
14'd471:data <=32'hFFE700B6;14'd472:data <=32'h000B00A9;14'd473:data <=32'h00270095;
14'd474:data <=32'h003D007D;14'd475:data <=32'h004D0062;14'd476:data <=32'h00540045;
14'd477:data <=32'h00530028;14'd478:data <=32'h004B000D;14'd479:data <=32'h003AFFF6;
14'd480:data <=32'h0023FFE7;14'd481:data <=32'h0009FFE1;14'd482:data <=32'hFFEEFFE6;
14'd483:data <=32'hFFD9FFF3;14'd484:data <=32'hFFC90007;14'd485:data <=32'hFFC3001D;
14'd486:data <=32'hFFC40034;14'd487:data <=32'hFFCD0047;14'd488:data <=32'hFFD90056;
14'd489:data <=32'hFFE50061;14'd490:data <=32'hFFF10069;14'd491:data <=32'hFFFE0070;
14'd492:data <=32'h000B0078;14'd493:data <=32'h001A007F;14'd494:data <=32'h002D0086;
14'd495:data <=32'h00450088;14'd496:data <=32'h005F0085;14'd497:data <=32'h0079007D;
14'd498:data <=32'h0093006E;14'd499:data <=32'h00AA0058;14'd500:data <=32'h00BB003E;
14'd501:data <=32'h00C80022;14'd502:data <=32'h00D00003;14'd503:data <=32'h00D3FFE2;
14'd504:data <=32'h00D0FFC0;14'd505:data <=32'h00C7FF9C;14'd506:data <=32'h00B6FF78;
14'd507:data <=32'h009AFF58;14'd508:data <=32'h0077FF3F;14'd509:data <=32'h004CFF32;
14'd510:data <=32'h0022FF31;14'd511:data <=32'hFFFAFF3E;14'd512:data <=32'h00B4FFB7;
14'd513:data <=32'h00B7FF81;14'd514:data <=32'h0097FF4B;14'd515:data <=32'hFFF4FF5C;
14'd516:data <=32'hFFCBFFA1;14'd517:data <=32'hFFD3FFB2;14'd518:data <=32'hFFDCFFBE;
14'd519:data <=32'hFFE7FFC1;14'd520:data <=32'hFFF0FFC0;14'd521:data <=32'hFFF8FFBB;
14'd522:data <=32'hFFFCFFB1;14'd523:data <=32'hFFFCFFA4;14'd524:data <=32'hFFF5FF93;
14'd525:data <=32'hFFE4FF83;14'd526:data <=32'hFFCBFF78;14'd527:data <=32'hFFADFF75;
14'd528:data <=32'hFF8BFF7E;14'd529:data <=32'hFF6BFF92;14'd530:data <=32'hFF54FFB1;
14'd531:data <=32'hFF48FFD6;14'd532:data <=32'hFF48FFFB;14'd533:data <=32'hFF50001E;
14'd534:data <=32'hFF62003A;14'd535:data <=32'hFF76004F;14'd536:data <=32'hFF8D005D;
14'd537:data <=32'hFFA30067;14'd538:data <=32'hFFB9006B;14'd539:data <=32'hFFCF006C;
14'd540:data <=32'hFFE40069;14'd541:data <=32'hFFF70063;14'd542:data <=32'h00080056;
14'd543:data <=32'h00140046;14'd544:data <=32'h00190033;14'd545:data <=32'h00190023;
14'd546:data <=32'h00140015;14'd547:data <=32'h000B000A;14'd548:data <=32'h00010004;
14'd549:data <=32'hFFF70001;14'd550:data <=32'hFFEFFFFE;14'd551:data <=32'hFFE6FFFD;
14'd552:data <=32'hFFDBFFFD;14'd553:data <=32'hFFCEFFFE;14'd554:data <=32'hFFBE0004;
14'd555:data <=32'hFFAD0010;14'd556:data <=32'hFF9C0024;14'd557:data <=32'hFF900040;
14'd558:data <=32'hFF8E0063;14'd559:data <=32'hFF970089;14'd560:data <=32'hFFAC00AC;
14'd561:data <=32'hFFCD00CC;14'd562:data <=32'hFFF600E2;14'd563:data <=32'h002500ED;
14'd564:data <=32'h005600EB;14'd565:data <=32'h008600DF;14'd566:data <=32'h00B300CA;
14'd567:data <=32'h00DB00A9;14'd568:data <=32'h00FD007E;14'd569:data <=32'h0115004B;
14'd570:data <=32'h01200014;14'd571:data <=32'h011DFFD9;14'd572:data <=32'h010BFFA1;
14'd573:data <=32'h00E8FF71;14'd574:data <=32'h00BCFF4F;14'd575:data <=32'h008BFF3C;
14'd576:data <=32'h008DFFDA;14'd577:data <=32'h0097FFC0;14'd578:data <=32'h00A2FF98;
14'd579:data <=32'h0086FF46;14'd580:data <=32'h0048FF76;14'd581:data <=32'h003AFF79;
14'd582:data <=32'h002DFF7C;14'd583:data <=32'h0023FF7D;14'd584:data <=32'h0018FF7E;
14'd585:data <=32'h000DFF81;14'd586:data <=32'h0005FF84;14'd587:data <=32'hFFFEFF87;
14'd588:data <=32'hFFF5FF86;14'd589:data <=32'hFFECFF85;14'd590:data <=32'hFFE0FF83;
14'd591:data <=32'hFFD0FF84;14'd592:data <=32'hFFBDFF8B;14'd593:data <=32'hFFAAFF97;
14'd594:data <=32'hFF9DFFA9;14'd595:data <=32'hFF96FFBF;14'd596:data <=32'hFF96FFD4;
14'd597:data <=32'hFF9DFFE5;14'd598:data <=32'hFFA8FFF1;14'd599:data <=32'hFFB2FFF6;
14'd600:data <=32'hFFBAFFF7;14'd601:data <=32'hFFBDFFF6;14'd602:data <=32'hFFBCFFF4;
14'd603:data <=32'hFFB9FFF6;14'd604:data <=32'hFFB7FFFC;14'd605:data <=32'hFFB60003;
14'd606:data <=32'hFFB6000A;14'd607:data <=32'hFFB80012;14'd608:data <=32'hFFBD0018;
14'd609:data <=32'hFFC2001D;14'd610:data <=32'hFFC70022;14'd611:data <=32'hFFCE0026;
14'd612:data <=32'hFFD6002A;14'd613:data <=32'hFFE0002A;14'd614:data <=32'hFFEA0028;
14'd615:data <=32'hFFF50020;14'd616:data <=32'hFFFA0012;14'd617:data <=32'hFFFB0001;
14'd618:data <=32'hFFF2FFF0;14'd619:data <=32'hFFDFFFE2;14'd620:data <=32'hFFC7FFDC;
14'd621:data <=32'hFFAAFFE0;14'd622:data <=32'hFF8DFFF0;14'd623:data <=32'hFF76000C;
14'd624:data <=32'hFF68002E;14'd625:data <=32'hFF660056;14'd626:data <=32'hFF6E007C;
14'd627:data <=32'hFF8200A1;14'd628:data <=32'hFF9E00C0;14'd629:data <=32'hFFBE00D9;
14'd630:data <=32'hFFE600E9;14'd631:data <=32'h001000F2;14'd632:data <=32'h003E00F2;
14'd633:data <=32'h006C00E8;14'd634:data <=32'h009600D2;14'd635:data <=32'h00BA00B2;
14'd636:data <=32'h00D4008A;14'd637:data <=32'h00E2005E;14'd638:data <=32'h00E40035;
14'd639:data <=32'h00DD0011;14'd640:data <=32'h00D20000;14'd641:data <=32'h00D4FFE2;
14'd642:data <=32'h00D7FFD5;14'd643:data <=32'h00F30012;14'd644:data <=32'h00D40023;
14'd645:data <=32'h00DF0006;14'd646:data <=32'h00E5FFE2;14'd647:data <=32'h00E3FFBA;
14'd648:data <=32'h00D5FF93;14'd649:data <=32'h00BFFF71;14'd650:data <=32'h00A1FF55;
14'd651:data <=32'h0080FF40;14'd652:data <=32'h005CFF32;14'd653:data <=32'h0036FF2A;
14'd654:data <=32'h000FFF2A;14'd655:data <=32'hFFE9FF32;14'd656:data <=32'hFFC4FF43;
14'd657:data <=32'hFFA4FF5D;14'd658:data <=32'hFF8EFF7F;14'd659:data <=32'hFF82FFA6;
14'd660:data <=32'hFF85FFCD;14'd661:data <=32'hFF92FFED;14'd662:data <=32'hFFAA0006;
14'd663:data <=32'hFFC50010;14'd664:data <=32'hFFDE0011;14'd665:data <=32'hFFF20009;
14'd666:data <=32'hFFFFFFFA;14'd667:data <=32'h0006FFEB;14'd668:data <=32'h0004FFDD;
14'd669:data <=32'hFFFEFFD1;14'd670:data <=32'hFFF7FFC8;14'd671:data <=32'hFFECFFC2;
14'd672:data <=32'hFFE2FFBF;14'd673:data <=32'hFFD4FFBF;14'd674:data <=32'hFFC8FFC4;
14'd675:data <=32'hFFBCFFCB;14'd676:data <=32'hFFB4FFD5;14'd677:data <=32'hFFAFFFE2;
14'd678:data <=32'hFFB0FFF0;14'd679:data <=32'hFFB5FFFA;14'd680:data <=32'hFFBD0000;
14'd681:data <=32'hFFC50000;14'd682:data <=32'hFFC9FFFC;14'd683:data <=32'hFFC9FFF4;
14'd684:data <=32'hFFC2FFEE;14'd685:data <=32'hFFB5FFEC;14'd686:data <=32'hFFA7FFEF;
14'd687:data <=32'hFF99FFFA;14'd688:data <=32'hFF8E0009;14'd689:data <=32'hFF88001D;
14'd690:data <=32'hFF890030;14'd691:data <=32'hFF8D0043;14'd692:data <=32'hFF950052;
14'd693:data <=32'hFF9D0060;14'd694:data <=32'hFFA7006C;14'd695:data <=32'hFFB10078;
14'd696:data <=32'hFFBC0083;14'd697:data <=32'hFFCA008F;14'd698:data <=32'hFFDA0097;
14'd699:data <=32'hFFEC009D;14'd700:data <=32'hFFFE009F;14'd701:data <=32'h000E009F;
14'd702:data <=32'h001C00A0;14'd703:data <=32'h002900A3;14'd704:data <=32'h00A300AC;
14'd705:data <=32'h00BF0096;14'd706:data <=32'h00C00081;14'd707:data <=32'h004F00BA;
14'd708:data <=32'h005000EA;14'd709:data <=32'h008300E5;14'd710:data <=32'h00B600D1;
14'd711:data <=32'h00E600AD;14'd712:data <=32'h0108007D;14'd713:data <=32'h011C0047;
14'd714:data <=32'h0123000F;14'd715:data <=32'h011DFFD7;14'd716:data <=32'h010CFFA3;
14'd717:data <=32'h00F1FF75;14'd718:data <=32'h00CBFF4D;14'd719:data <=32'h009EFF30;
14'd720:data <=32'h006AFF1C;14'd721:data <=32'h0035FF1B;14'd722:data <=32'h0000FF26;
14'd723:data <=32'hFFD5FF40;14'd724:data <=32'hFFB5FF63;14'd725:data <=32'hFFA4FF8C;
14'd726:data <=32'hFFA1FFB1;14'd727:data <=32'hFFA9FFD2;14'd728:data <=32'hFFB8FFE9;
14'd729:data <=32'hFFCAFFF8;14'd730:data <=32'hFFDB0000;14'd731:data <=32'hFFEA0002;
14'd732:data <=32'hFFF80003;14'd733:data <=32'h00030000;14'd734:data <=32'h000EFFFB;
14'd735:data <=32'h0018FFF3;14'd736:data <=32'h001FFFE9;14'd737:data <=32'h0024FFDC;
14'd738:data <=32'h0025FFCE;14'd739:data <=32'h0020FFBE;14'd740:data <=32'h0018FFB2;
14'd741:data <=32'h000CFFA8;14'd742:data <=32'h0000FFA1;14'd743:data <=32'hFFF3FF9D;
14'd744:data <=32'hFFE5FF99;14'd745:data <=32'hFFD8FF97;14'd746:data <=32'hFFC8FF94;
14'd747:data <=32'hFFB6FF95;14'd748:data <=32'hFFA1FF99;14'd749:data <=32'hFF8CFFA3;
14'd750:data <=32'hFF75FFB5;14'd751:data <=32'hFF64FFCD;14'd752:data <=32'hFF5BFFEB;
14'd753:data <=32'hFF5B000B;14'd754:data <=32'hFF640027;14'd755:data <=32'hFF750040;
14'd756:data <=32'hFF8B004F;14'd757:data <=32'hFFA10056;14'd758:data <=32'hFFB40056;
14'd759:data <=32'hFFC30051;14'd760:data <=32'hFFCB004A;14'd761:data <=32'hFFD00043;
14'd762:data <=32'hFFD1003D;14'd763:data <=32'hFFCE0038;14'd764:data <=32'hFFC80035;
14'd765:data <=32'hFFBD0037;14'd766:data <=32'hFFB1003D;14'd767:data <=32'hFFA5004D;
14'd768:data <=32'hFFCE00AB;14'd769:data <=32'hFFE000C0;14'd770:data <=32'hFFF200BB;
14'd771:data <=32'hFFC10079;14'd772:data <=32'hFFAA00C1;14'd773:data <=32'hFFCE00DD;
14'd774:data <=32'hFFFB00EE;14'd775:data <=32'h002C00F1;14'd776:data <=32'h005A00E6;
14'd777:data <=32'h008400D1;14'd778:data <=32'h00A500B5;14'd779:data <=32'h00BF0094;
14'd780:data <=32'h00D3006F;14'd781:data <=32'h00DE0048;14'd782:data <=32'h00E2001F;
14'd783:data <=32'h00DDFFF6;14'd784:data <=32'h00CFFFD0;14'd785:data <=32'h00B8FFAF;
14'd786:data <=32'h009BFF98;14'd787:data <=32'h007AFF8B;14'd788:data <=32'h005CFF87;
14'd789:data <=32'h0042FF89;14'd790:data <=32'h002EFF90;14'd791:data <=32'h0020FF99;
14'd792:data <=32'h0015FF9F;14'd793:data <=32'h000BFFA5;14'd794:data <=32'hFFFFFFAB;
14'd795:data <=32'hFFF4FFB2;14'd796:data <=32'hFFEAFFBD;14'd797:data <=32'hFFE1FFCC;
14'd798:data <=32'hFFDEFFDE;14'd799:data <=32'hFFE2FFF1;14'd800:data <=32'hFFEC0001;
14'd801:data <=32'hFFFA000C;14'd802:data <=32'h000E0012;14'd803:data <=32'h00210011;
14'd804:data <=32'h00340009;14'd805:data <=32'h0043FFFC;14'd806:data <=32'h0051FFEB;
14'd807:data <=32'h0059FFD5;14'd808:data <=32'h005CFFBD;14'd809:data <=32'h005AFFA1;
14'd810:data <=32'h0051FF84;14'd811:data <=32'h003DFF69;14'd812:data <=32'h0020FF51;
14'd813:data <=32'hFFFCFF41;14'd814:data <=32'hFFD1FF3C;14'd815:data <=32'hFFA6FF46;
14'd816:data <=32'hFF80FF5B;14'd817:data <=32'hFF62FF7A;14'd818:data <=32'hFF4FFF9E;
14'd819:data <=32'hFF49FFC5;14'd820:data <=32'hFF4DFFE7;14'd821:data <=32'hFF590003;
14'd822:data <=32'hFF670017;14'd823:data <=32'hFF770024;14'd824:data <=32'hFF86002D;
14'd825:data <=32'hFF940032;14'd826:data <=32'hFF9E0034;14'd827:data <=32'hFFA70033;
14'd828:data <=32'hFFAC0030;14'd829:data <=32'hFFAD002D;14'd830:data <=32'hFFA9002A;
14'd831:data <=32'hFFA0002D;14'd832:data <=32'hFFA60002;14'd833:data <=32'hFF860011;
14'd834:data <=32'hFF7F002D;14'd835:data <=32'hFFB4005F;14'd836:data <=32'hFF950098;
14'd837:data <=32'hFFAE00AC;14'd838:data <=32'hFFCE00B6;14'd839:data <=32'hFFEF00B9;
14'd840:data <=32'h000E00B1;14'd841:data <=32'h002600A3;14'd842:data <=32'h00370092;
14'd843:data <=32'h00420081;14'd844:data <=32'h00490073;14'd845:data <=32'h004E0067;
14'd846:data <=32'h0053005C;14'd847:data <=32'h00570052;14'd848:data <=32'h005B0048;
14'd849:data <=32'h005D003D;14'd850:data <=32'h005D0036;14'd851:data <=32'h005D002F;
14'd852:data <=32'h005E002A;14'd853:data <=32'h00620027;14'd854:data <=32'h006B0020;
14'd855:data <=32'h00740017;14'd856:data <=32'h007D0006;14'd857:data <=32'h0080FFF0;
14'd858:data <=32'h007CFFD8;14'd859:data <=32'h006FFFC0;14'd860:data <=32'h005BFFAE;
14'd861:data <=32'h0041FFA4;14'd862:data <=32'h0026FFA3;14'd863:data <=32'h000CFFAC;
14'd864:data <=32'hFFFAFFBC;14'd865:data <=32'hFFEFFFD0;14'd866:data <=32'hFFECFFE5;
14'd867:data <=32'hFFEFFFF9;14'd868:data <=32'hFFF9000A;14'd869:data <=32'h00080017;
14'd870:data <=32'h001B001F;14'd871:data <=32'h002F0021;14'd872:data <=32'h0047001E;
14'd873:data <=32'h005D0011;14'd874:data <=32'h0071FFFD;14'd875:data <=32'h007EFFE2;
14'd876:data <=32'h0084FFC1;14'd877:data <=32'h007EFFA0;14'd878:data <=32'h006DFF7F;
14'd879:data <=32'h0055FF66;14'd880:data <=32'h0038FF56;14'd881:data <=32'h0018FF4F;
14'd882:data <=32'hFFFCFF4F;14'd883:data <=32'hFFE3FF54;14'd884:data <=32'hFFCEFF5B;
14'd885:data <=32'hFFBDFF63;14'd886:data <=32'hFFACFF6A;14'd887:data <=32'hFF9BFF71;
14'd888:data <=32'hFF87FF79;14'd889:data <=32'hFF73FF85;14'd890:data <=32'hFF61FF96;
14'd891:data <=32'hFF50FFAB;14'd892:data <=32'hFF44FFC2;14'd893:data <=32'hFF3CFFDC;
14'd894:data <=32'hFF37FFF5;14'd895:data <=32'hFF34000F;14'd896:data <=32'hFFEBFFE2;
14'd897:data <=32'hFFCBFFCC;14'd898:data <=32'hFF9DFFD0;14'd899:data <=32'hFF3B004D;
14'd900:data <=32'hFF26009A;14'd901:data <=32'hFF4E00BD;14'd902:data <=32'hFF7F00D4;
14'd903:data <=32'hFFB300DD;14'd904:data <=32'hFFE300D5;14'd905:data <=32'h000C00C0;
14'd906:data <=32'h002900A2;14'd907:data <=32'h00380083;14'd908:data <=32'h003E0067;
14'd909:data <=32'h003B004F;14'd910:data <=32'h0033003C;14'd911:data <=32'h0028002F;
14'd912:data <=32'h001D0028;14'd913:data <=32'h00110026;14'd914:data <=32'h00060029;
14'd915:data <=32'hFFFD0031;14'd916:data <=32'hFFFA003F;14'd917:data <=32'hFFFC004E;
14'd918:data <=32'h0007005E;14'd919:data <=32'h001A0069;14'd920:data <=32'h0032006D;
14'd921:data <=32'h004B0066;14'd922:data <=32'h00610056;14'd923:data <=32'h006F0040;
14'd924:data <=32'h00760026;14'd925:data <=32'h0072000F;14'd926:data <=32'h0069FFFA;
14'd927:data <=32'h005CFFEC;14'd928:data <=32'h004CFFE5;14'd929:data <=32'h003FFFE3;
14'd930:data <=32'h0035FFE2;14'd931:data <=32'h002BFFE6;14'd932:data <=32'h0024FFE9;
14'd933:data <=32'h001FFFEE;14'd934:data <=32'h001BFFF5;14'd935:data <=32'h001AFFFD;
14'd936:data <=32'h001D0005;14'd937:data <=32'h0022000D;14'd938:data <=32'h002C0012;
14'd939:data <=32'h00390012;14'd940:data <=32'h00450010;14'd941:data <=32'h00500008;
14'd942:data <=32'h0059FFFD;14'd943:data <=32'h005FFFF2;14'd944:data <=32'h0063FFE8;
14'd945:data <=32'h0067FFDE;14'd946:data <=32'h006AFFD4;14'd947:data <=32'h0072FFC6;
14'd948:data <=32'h007AFFB5;14'd949:data <=32'h007EFF9D;14'd950:data <=32'h007EFF7E;
14'd951:data <=32'h0074FF5A;14'd952:data <=32'h005EFF37;14'd953:data <=32'h003CFF18;
14'd954:data <=32'h0012FF01;14'd955:data <=32'hFFE1FEF6;14'd956:data <=32'hFFADFEF6;
14'd957:data <=32'hFF7AFF02;14'd958:data <=32'hFF4AFF1A;14'd959:data <=32'hFF1FFF3B;
14'd960:data <=32'hFFC6FFC6;14'd961:data <=32'hFFB5FFB1;14'd962:data <=32'hFF92FF95;
14'd963:data <=32'hFF07FF74;14'd964:data <=32'hFEC9FFD4;14'd965:data <=32'hFED20015;
14'd966:data <=32'hFEEA004F;14'd967:data <=32'hFF10007E;14'd968:data <=32'hFF3F009E;
14'd969:data <=32'hFF6E00AD;14'd970:data <=32'hFF9A00AE;14'd971:data <=32'hFFBF00A5;
14'd972:data <=32'hFFDB0097;14'd973:data <=32'hFFEF0088;14'd974:data <=32'hFFFE0077;
14'd975:data <=32'h00080068;14'd976:data <=32'h000E0059;14'd977:data <=32'h0010004B;
14'd978:data <=32'h000E003E;14'd979:data <=32'h00080035;14'd980:data <=32'h00010031;
14'd981:data <=32'hFFF90033;14'd982:data <=32'hFFF60039;14'd983:data <=32'hFFF60040;
14'd984:data <=32'hFFFD0048;14'd985:data <=32'h0006004B;14'd986:data <=32'h0011004A;
14'd987:data <=32'h001A0044;14'd988:data <=32'h001D003D;14'd989:data <=32'h001D0037;
14'd990:data <=32'h001C0033;14'd991:data <=32'h00190033;14'd992:data <=32'h00190037;
14'd993:data <=32'h001C003C;14'd994:data <=32'h00240040;14'd995:data <=32'h002E0040;
14'd996:data <=32'h003A003D;14'd997:data <=32'h00440036;14'd998:data <=32'h004B002C;
14'd999:data <=32'h004E0020;14'd1000:data <=32'h004D0016;14'd1001:data <=32'h004B000D;
14'd1002:data <=32'h00470005;14'd1003:data <=32'h00430000;14'd1004:data <=32'h003DFFFD;
14'd1005:data <=32'h0037FFFB;14'd1006:data <=32'h0031FFFB;14'd1007:data <=32'h002A0000;
14'd1008:data <=32'h00270009;14'd1009:data <=32'h00280016;14'd1010:data <=32'h00320023;
14'd1011:data <=32'h0044002F;14'd1012:data <=32'h005E0035;14'd1013:data <=32'h007D002F;
14'd1014:data <=32'h009F001D;14'd1015:data <=32'h00BAFFFD;14'd1016:data <=32'h00CCFFD3;
14'd1017:data <=32'h00D2FFA2;14'd1018:data <=32'h00C7FF6F;14'd1019:data <=32'h00B0FF40;
14'd1020:data <=32'h008EFF18;14'd1021:data <=32'h0063FEF9;14'd1022:data <=32'h0031FEE3;
14'd1023:data <=32'hFFFBFED8;14'd1024:data <=32'h0012FF3F;14'd1025:data <=32'hFFF0FF1F;
14'd1026:data <=32'hFFD7FF08;14'd1027:data <=32'hFFD6FEF1;14'd1028:data <=32'hFF7AFF27;
14'd1029:data <=32'hFF5AFF48;14'd1030:data <=32'hFF47FF6E;14'd1031:data <=32'hFF3EFF95;
14'd1032:data <=32'hFF3EFFB6;14'd1033:data <=32'hFF43FFD1;14'd1034:data <=32'hFF4AFFE6;
14'd1035:data <=32'hFF4FFFF8;14'd1036:data <=32'hFF520009;14'd1037:data <=32'hFF56001B;
14'd1038:data <=32'hFF5C0031;14'd1039:data <=32'hFF660046;14'd1040:data <=32'hFF74005A;
14'd1041:data <=32'hFF88006B;14'd1042:data <=32'hFF9E0075;14'd1043:data <=32'hFFB5007B;
14'd1044:data <=32'hFFCB007C;14'd1045:data <=32'hFFDF007B;14'd1046:data <=32'hFFF10076;
14'd1047:data <=32'h0003006E;14'd1048:data <=32'h00130063;14'd1049:data <=32'h00220054;
14'd1050:data <=32'h002C0041;14'd1051:data <=32'h002E002A;14'd1052:data <=32'h00280015;
14'd1053:data <=32'h001A0002;14'd1054:data <=32'h0006FFF8;14'd1055:data <=32'hFFF0FFF8;
14'd1056:data <=32'hFFDB0001;14'd1057:data <=32'hFFCC0012;14'd1058:data <=32'hFFC50028;
14'd1059:data <=32'hFFC7003F;14'd1060:data <=32'hFFD10052;14'd1061:data <=32'hFFE10061;
14'd1062:data <=32'hFFF3006A;14'd1063:data <=32'h0006006E;14'd1064:data <=32'h0018006C;
14'd1065:data <=32'h00280067;14'd1066:data <=32'h00360060;14'd1067:data <=32'h00420056;
14'd1068:data <=32'h004B004A;14'd1069:data <=32'h0050003C;14'd1070:data <=32'h00500030;
14'd1071:data <=32'h004E0025;14'd1072:data <=32'h00460020;14'd1073:data <=32'h003F001F;
14'd1074:data <=32'h003B0024;14'd1075:data <=32'h003D002F;14'd1076:data <=32'h00470038;
14'd1077:data <=32'h0059003F;14'd1078:data <=32'h0070003E;14'd1079:data <=32'h00880034;
14'd1080:data <=32'h009E001F;14'd1081:data <=32'h00AE0004;14'd1082:data <=32'h00B6FFE3;
14'd1083:data <=32'h00B4FFC3;14'd1084:data <=32'h00ACFFA4;14'd1085:data <=32'h009FFF89;
14'd1086:data <=32'h008DFF71;14'd1087:data <=32'h0078FF5D;14'd1088:data <=32'h00E0FF76;
14'd1089:data <=32'h00D3FF31;14'd1090:data <=32'h00B0FF08;14'd1091:data <=32'h0066FF5F;
14'd1092:data <=32'h0021FF78;14'd1093:data <=32'h0017FF7B;14'd1094:data <=32'h0010FF7D;
14'd1095:data <=32'h0009FF7D;14'd1096:data <=32'h0005FF79;14'd1097:data <=32'hFFFEFF6F;
14'd1098:data <=32'hFFF3FF62;14'd1099:data <=32'hFFDDFF56;14'd1100:data <=32'hFFC1FF4E;
14'd1101:data <=32'hFF9CFF4F;14'd1102:data <=32'hFF78FF5C;14'd1103:data <=32'hFF56FF74;
14'd1104:data <=32'hFF3CFF97;14'd1105:data <=32'hFF2DFFBE;14'd1106:data <=32'hFF28FFE9;
14'd1107:data <=32'hFF2D0011;14'd1108:data <=32'hFF3B0037;14'd1109:data <=32'hFF4F0057;
14'd1110:data <=32'hFF6B0072;14'd1111:data <=32'hFF8B0087;14'd1112:data <=32'hFFAF0091;
14'd1113:data <=32'hFFD60093;14'd1114:data <=32'hFFFB0088;14'd1115:data <=32'h001A0072;
14'd1116:data <=32'h002F0056;14'd1117:data <=32'h00380034;14'd1118:data <=32'h00360015;
14'd1119:data <=32'h0027FFF9;14'd1120:data <=32'h0012FFE7;14'd1121:data <=32'hFFF9FFDF;
14'd1122:data <=32'hFFE2FFE1;14'd1123:data <=32'hFFCFFFE9;14'd1124:data <=32'hFFC0FFF5;
14'd1125:data <=32'hFFB70003;14'd1126:data <=32'hFFB00012;14'd1127:data <=32'hFFAD0022;
14'd1128:data <=32'hFFAB0031;14'd1129:data <=32'hFFAC0041;14'd1130:data <=32'hFFB00054;
14'd1131:data <=32'hFFB90065;14'd1132:data <=32'hFFC50074;14'd1133:data <=32'hFFD50082;
14'd1134:data <=32'hFFE8008C;14'd1135:data <=32'hFFFA0091;14'd1136:data <=32'h000D0095;
14'd1137:data <=32'h00200097;14'd1138:data <=32'h00320098;14'd1139:data <=32'h00470097;
14'd1140:data <=32'h005F0095;14'd1141:data <=32'h007A008D;14'd1142:data <=32'h0096007E;
14'd1143:data <=32'h00AF0065;14'd1144:data <=32'h00C30046;14'd1145:data <=32'h00CC0020;
14'd1146:data <=32'h00CCFFFA;14'd1147:data <=32'h00C1FFD6;14'd1148:data <=32'h00ADFFBA;
14'd1149:data <=32'h0095FFA5;14'd1150:data <=32'h007CFF9B;14'd1151:data <=32'h0066FF96;
14'd1152:data <=32'h00E0003A;14'd1153:data <=32'h01060004;14'd1154:data <=32'h0105FFC1;
14'd1155:data <=32'h0065FF95;14'd1156:data <=32'h0024FFBA;14'd1157:data <=32'h0024FFC8;
14'd1158:data <=32'h002BFFD3;14'd1159:data <=32'h0037FFD9;14'd1160:data <=32'h0048FFD7;
14'd1161:data <=32'h005AFFCB;14'd1162:data <=32'h0066FFB3;14'd1163:data <=32'h0068FF95;
14'd1164:data <=32'h005EFF73;14'd1165:data <=32'h0046FF55;14'd1166:data <=32'h0025FF3E;
14'd1167:data <=32'hFFFDFF34;14'd1168:data <=32'hFFD4FF36;14'd1169:data <=32'hFFAEFF42;
14'd1170:data <=32'hFF8EFF57;14'd1171:data <=32'hFF74FF71;14'd1172:data <=32'hFF61FF8F;
14'd1173:data <=32'hFF54FFAF;14'd1174:data <=32'hFF4FFFD1;14'd1175:data <=32'hFF51FFF4;
14'd1176:data <=32'hFF5B0015;14'd1177:data <=32'hFF6F0032;14'd1178:data <=32'hFF880047;
14'd1179:data <=32'hFFA60054;14'd1180:data <=32'hFFC20055;14'd1181:data <=32'hFFDC004F;
14'd1182:data <=32'hFFF00042;14'd1183:data <=32'hFFFC0033;14'd1184:data <=32'h00020023;
14'd1185:data <=32'h00030016;14'd1186:data <=32'h0002000C;14'd1187:data <=32'h00010003;
14'd1188:data <=32'hFFFFFFFA;14'd1189:data <=32'hFFFCFFEF;14'd1190:data <=32'hFFF4FFE4;
14'd1191:data <=32'hFFE9FFD8;14'd1192:data <=32'hFFD8FFCF;14'd1193:data <=32'hFFC2FFCB;
14'd1194:data <=32'hFFA9FFCF;14'd1195:data <=32'hFF8FFFDB;14'd1196:data <=32'hFF79FFEF;
14'd1197:data <=32'hFF69000A;14'd1198:data <=32'hFF5E002A;14'd1199:data <=32'hFF5B004B;
14'd1200:data <=32'hFF5F0070;14'd1201:data <=32'hFF6B0094;14'd1202:data <=32'hFF8100B8;
14'd1203:data <=32'hFF9E00D9;14'd1204:data <=32'hFFC500F4;14'd1205:data <=32'hFFF40106;
14'd1206:data <=32'h002B010D;14'd1207:data <=32'h00630103;14'd1208:data <=32'h009700EB;
14'd1209:data <=32'h00C400C3;14'd1210:data <=32'h00E10093;14'd1211:data <=32'h00F0005D;
14'd1212:data <=32'h00EF002A;14'd1213:data <=32'h00E0FFFE;14'd1214:data <=32'h00CAFFDC;
14'd1215:data <=32'h00B0FFC3;14'd1216:data <=32'h007B0056;14'd1217:data <=32'h009D004B;
14'd1218:data <=32'h00C10026;14'd1219:data <=32'h00C0FFBD;14'd1220:data <=32'h0077FFCD;
14'd1221:data <=32'h006AFFCB;14'd1222:data <=32'h0060FFCD;14'd1223:data <=32'h005BFFD1;
14'd1224:data <=32'h005CFFD3;14'd1225:data <=32'h0062FFD1;14'd1226:data <=32'h0068FFC8;
14'd1227:data <=32'h006CFFB7;14'd1228:data <=32'h0069FFA3;14'd1229:data <=32'h005EFF8F;
14'd1230:data <=32'h004BFF7D;14'd1231:data <=32'h0033FF73;14'd1232:data <=32'h001BFF71;
14'd1233:data <=32'h0005FF74;14'd1234:data <=32'hFFF4FF7C;14'd1235:data <=32'hFFE6FF87;
14'd1236:data <=32'hFFDCFF90;14'd1237:data <=32'hFFD3FF99;14'd1238:data <=32'hFFCBFFA1;
14'd1239:data <=32'hFFC3FFAB;14'd1240:data <=32'hFFBEFFB6;14'd1241:data <=32'hFFB8FFC1;
14'd1242:data <=32'hFFB8FFCC;14'd1243:data <=32'hFFB9FFD7;14'd1244:data <=32'hFFBCFFDD;
14'd1245:data <=32'hFFBEFFE2;14'd1246:data <=32'hFFC0FFE5;14'd1247:data <=32'hFFBEFFEA;
14'd1248:data <=32'hFFBBFFF0;14'd1249:data <=32'hFFBBFFFA;14'd1250:data <=32'hFFBF0006;
14'd1251:data <=32'hFFC60010;14'd1252:data <=32'hFFD40019;14'd1253:data <=32'hFFE50019;
14'd1254:data <=32'hFFF70014;14'd1255:data <=32'h00050005;14'd1256:data <=32'h000CFFF0;
14'd1257:data <=32'h000AFFD9;14'd1258:data <=32'hFFFFFFC2;14'd1259:data <=32'hFFEBFFB0;
14'd1260:data <=32'hFFCFFFA5;14'd1261:data <=32'hFFB1FFA2;14'd1262:data <=32'hFF92FFA8;
14'd1263:data <=32'hFF73FFB7;14'd1264:data <=32'hFF58FFCE;14'd1265:data <=32'hFF41FFEC;
14'd1266:data <=32'hFF300012;14'd1267:data <=32'hFF28003D;14'd1268:data <=32'hFF2C006D;
14'd1269:data <=32'hFF3C009D;14'd1270:data <=32'hFF5B00C8;14'd1271:data <=32'hFF8400EA;
14'd1272:data <=32'hFFB500FF;14'd1273:data <=32'hFFE90105;14'd1274:data <=32'h001A00FE;
14'd1275:data <=32'h004400EB;14'd1276:data <=32'h006400D3;14'd1277:data <=32'h007C00B8;
14'd1278:data <=32'h008B009F;14'd1279:data <=32'h00960086;14'd1280:data <=32'h0087006A;
14'd1281:data <=32'h0099005D;14'd1282:data <=32'h00AC0059;14'd1283:data <=32'h00C4008F;
14'd1284:data <=32'h00A0008F;14'd1285:data <=32'h00B30077;14'd1286:data <=32'h00C2005D;
14'd1287:data <=32'h00CD0041;14'd1288:data <=32'h00D50023;14'd1289:data <=32'h00D80004;
14'd1290:data <=32'h00D9FFE1;14'd1291:data <=32'h00D1FFBD;14'd1292:data <=32'h00BFFF99;
14'd1293:data <=32'h00A4FF78;14'd1294:data <=32'h007FFF62;14'd1295:data <=32'h0055FF56;
14'd1296:data <=32'h002DFF58;14'd1297:data <=32'h0009FF66;14'd1298:data <=32'hFFEEFF7C;
14'd1299:data <=32'hFFDFFF96;14'd1300:data <=32'hFFD9FFAF;14'd1301:data <=32'hFFDCFFC5;
14'd1302:data <=32'hFFE3FFD5;14'd1303:data <=32'hFFECFFE1;14'd1304:data <=32'hFFF7FFE6;
14'd1305:data <=32'h0002FFE8;14'd1306:data <=32'h000CFFE7;14'd1307:data <=32'h0016FFE0;
14'd1308:data <=32'h001CFFD7;14'd1309:data <=32'h001EFFCA;14'd1310:data <=32'h001AFFBB;
14'd1311:data <=32'h0010FFB0;14'd1312:data <=32'h0000FFA7;14'd1313:data <=32'hFFEDFFA6;
14'd1314:data <=32'hFFDCFFAC;14'd1315:data <=32'hFFCFFFB7;14'd1316:data <=32'hFFC9FFC7;
14'd1317:data <=32'hFFC9FFD6;14'd1318:data <=32'hFFD0FFE3;14'd1319:data <=32'hFFDBFFE7;
14'd1320:data <=32'hFFE6FFE6;14'd1321:data <=32'hFFEDFFDF;14'd1322:data <=32'hFFEFFFD4;
14'd1323:data <=32'hFFEDFFC9;14'd1324:data <=32'hFFE5FFC0;14'd1325:data <=32'hFFDAFFB8;
14'd1326:data <=32'hFFCCFFB5;14'd1327:data <=32'hFFBDFFB3;14'd1328:data <=32'hFFAEFFB4;
14'd1329:data <=32'hFF9DFFB9;14'd1330:data <=32'hFF8BFFC2;14'd1331:data <=32'hFF79FFCF;
14'd1332:data <=32'hFF69FFE2;14'd1333:data <=32'hFF5FFFF8;14'd1334:data <=32'hFF5A0013;
14'd1335:data <=32'hFF5C002E;14'd1336:data <=32'hFF640046;14'd1337:data <=32'hFF710059;
14'd1338:data <=32'hFF7D0068;14'd1339:data <=32'hFF880073;14'd1340:data <=32'hFF91007D;
14'd1341:data <=32'hFF97008B;14'd1342:data <=32'hFF9E009C;14'd1343:data <=32'hFFAA00B0;
14'd1344:data <=32'h002700D3;14'd1345:data <=32'h004600D1;14'd1346:data <=32'h004F00C6;
14'd1347:data <=32'hFFDB00E3;14'd1348:data <=32'hFFCD010B;14'd1349:data <=32'hFFFF0118;
14'd1350:data <=32'h0033011A;14'd1351:data <=32'h00670110;14'd1352:data <=32'h009900FB;
14'd1353:data <=32'h00C800DB;14'd1354:data <=32'h00EF00B1;14'd1355:data <=32'h010C007C;
14'd1356:data <=32'h011B0040;14'd1357:data <=32'h011A0001;14'd1358:data <=32'h0106FFC7;
14'd1359:data <=32'h00E3FF96;14'd1360:data <=32'h00B7FF74;14'd1361:data <=32'h0085FF63;
14'd1362:data <=32'h0057FF61;14'd1363:data <=32'h002EFF6B;14'd1364:data <=32'h000FFF7D;
14'd1365:data <=32'hFFF9FF92;14'd1366:data <=32'hFFECFFA9;14'd1367:data <=32'hFFE5FFBF;
14'd1368:data <=32'hFFE3FFD4;14'd1369:data <=32'hFFE7FFE6;14'd1370:data <=32'hFFF0FFF7;
14'd1371:data <=32'hFFFD0004;14'd1372:data <=32'h000D000A;14'd1373:data <=32'h001E000A;
14'd1374:data <=32'h002D0003;14'd1375:data <=32'h0039FFF7;14'd1376:data <=32'h003DFFEA;
14'd1377:data <=32'h003EFFDA;14'd1378:data <=32'h003AFFCF;14'd1379:data <=32'h0033FFC6;
14'd1380:data <=32'h002FFFC1;14'd1381:data <=32'h002BFFBD;14'd1382:data <=32'h0028FFB8;
14'd1383:data <=32'h0027FFB0;14'd1384:data <=32'h0023FFA5;14'd1385:data <=32'h001CFF98;
14'd1386:data <=32'h000EFF8C;14'd1387:data <=32'hFFFBFF83;14'd1388:data <=32'hFFE7FF80;
14'd1389:data <=32'hFFD0FF83;14'd1390:data <=32'hFFBCFF8C;14'd1391:data <=32'hFFABFF9A;
14'd1392:data <=32'hFFA1FFAA;14'd1393:data <=32'hFF9AFFBA;14'd1394:data <=32'hFF97FFC9;
14'd1395:data <=32'hFF96FFD7;14'd1396:data <=32'hFF99FFE2;14'd1397:data <=32'hFF9DFFED;
14'd1398:data <=32'hFFA2FFF5;14'd1399:data <=32'hFFA9FFFB;14'd1400:data <=32'hFFB0FFFB;
14'd1401:data <=32'hFFB5FFF6;14'd1402:data <=32'hFFB5FFEF;14'd1403:data <=32'hFFADFFE4;
14'd1404:data <=32'hFF9DFFDC;14'd1405:data <=32'hFF84FFDC;14'd1406:data <=32'hFF67FFE7;
14'd1407:data <=32'hFF4BFFFF;14'd1408:data <=32'hFF6C0075;14'd1409:data <=32'hFF710092;
14'd1410:data <=32'hFF820097;14'd1411:data <=32'hFF600049;14'd1412:data <=32'hFF310084;
14'd1413:data <=32'hFF4600AE;14'd1414:data <=32'hFF6500D3;14'd1415:data <=32'hFF8D00EF;
14'd1416:data <=32'hFFB90104;14'd1417:data <=32'hFFEB0110;14'd1418:data <=32'h001F010F;
14'd1419:data <=32'h00540102;14'd1420:data <=32'h008100E7;14'd1421:data <=32'h00A800C1;
14'd1422:data <=32'h00C00094;14'd1423:data <=32'h00CA0064;14'd1424:data <=32'h00C70039;
14'd1425:data <=32'h00BB0015;14'd1426:data <=32'h00A9FFFA;14'd1427:data <=32'h0096FFE6;
14'd1428:data <=32'h0084FFD8;14'd1429:data <=32'h0074FFCE;14'd1430:data <=32'h0064FFC6;
14'd1431:data <=32'h0054FFBE;14'd1432:data <=32'h0043FFBB;14'd1433:data <=32'h0031FFBA;
14'd1434:data <=32'h001FFFBE;14'd1435:data <=32'h0011FFC7;14'd1436:data <=32'h0006FFD3;
14'd1437:data <=32'h0000FFE1;14'd1438:data <=32'hFFFFFFEE;14'd1439:data <=32'h0000FFFA;
14'd1440:data <=32'h00050004;14'd1441:data <=32'h000C000D;14'd1442:data <=32'h00140015;
14'd1443:data <=32'h0020001C;14'd1444:data <=32'h002F0021;14'd1445:data <=32'h00420022;
14'd1446:data <=32'h0058001C;14'd1447:data <=32'h006F000D;14'd1448:data <=32'h0080FFF6;
14'd1449:data <=32'h008BFFD7;14'd1450:data <=32'h008CFFB4;14'd1451:data <=32'h0082FF90;
14'd1452:data <=32'h006CFF71;14'd1453:data <=32'h004FFF5A;14'd1454:data <=32'h002CFF4D;
14'd1455:data <=32'h0008FF49;14'd1456:data <=32'hFFE8FF50;14'd1457:data <=32'hFFCBFF5D;
14'd1458:data <=32'hFFB5FF6E;14'd1459:data <=32'hFFA4FF81;14'd1460:data <=32'hFF99FF96;
14'd1461:data <=32'hFF94FFAC;14'd1462:data <=32'hFF94FFC1;14'd1463:data <=32'hFF99FFD3;
14'd1464:data <=32'hFFA4FFE0;14'd1465:data <=32'hFFB1FFE5;14'd1466:data <=32'hFFBDFFE2;
14'd1467:data <=32'hFFC4FFD9;14'd1468:data <=32'hFFC3FFCA;14'd1469:data <=32'hFFB6FFBC;
14'd1470:data <=32'hFFA0FFB4;14'd1471:data <=32'hFF85FFB6;14'd1472:data <=32'hFF98FFAE;
14'd1473:data <=32'hFF6EFFB4;14'd1474:data <=32'hFF5DFFCC;14'd1475:data <=32'hFF820000;
14'd1476:data <=32'hFF490029;14'd1477:data <=32'hFF530044;14'd1478:data <=32'hFF61005B;
14'd1479:data <=32'hFF72006E;14'd1480:data <=32'hFF84007F;14'd1481:data <=32'hFF97008C;
14'd1482:data <=32'hFFAD0097;14'd1483:data <=32'hFFC6009D;14'd1484:data <=32'hFFDE009E;
14'd1485:data <=32'hFFF40099;14'd1486:data <=32'h0007008F;14'd1487:data <=32'h00130084;
14'd1488:data <=32'h001A007A;14'd1489:data <=32'h001E0073;14'd1490:data <=32'h00220071;
14'd1491:data <=32'h002A0073;14'd1492:data <=32'h00380074;14'd1493:data <=32'h00480071;
14'd1494:data <=32'h005C0068;14'd1495:data <=32'h006E0058;14'd1496:data <=32'h007B0041;
14'd1497:data <=32'h00800028;14'd1498:data <=32'h007E000E;14'd1499:data <=32'h0075FFF7;
14'd1500:data <=32'h0066FFE5;14'd1501:data <=32'h0054FFD8;14'd1502:data <=32'h0041FFCF;
14'd1503:data <=32'h002DFFCD;14'd1504:data <=32'h0018FFCF;14'd1505:data <=32'h0006FFD8;
14'd1506:data <=32'hFFF7FFE6;14'd1507:data <=32'hFFECFFFA;14'd1508:data <=32'hFFEB0014;
14'd1509:data <=32'hFFF2002D;14'd1510:data <=32'h00030042;14'd1511:data <=32'h001D0052;
14'd1512:data <=32'h003D0057;14'd1513:data <=32'h005E0051;14'd1514:data <=32'h007B003F;
14'd1515:data <=32'h00920025;14'd1516:data <=32'h009F0005;14'd1517:data <=32'h00A2FFE5;
14'd1518:data <=32'h009DFFC7;14'd1519:data <=32'h0092FFAC;14'd1520:data <=32'h0083FF96;
14'd1521:data <=32'h0072FF84;14'd1522:data <=32'h0062FF75;14'd1523:data <=32'h004EFF6A;
14'd1524:data <=32'h003AFF5F;14'd1525:data <=32'h0024FF5A;14'd1526:data <=32'h000EFF57;
14'd1527:data <=32'hFFF8FF59;14'd1528:data <=32'hFFE6FF5D;14'd1529:data <=32'hFFD6FF62;
14'd1530:data <=32'hFFC9FF67;14'd1531:data <=32'hFFBBFF6A;14'd1532:data <=32'hFFABFF6C;
14'd1533:data <=32'hFF98FF6F;14'd1534:data <=32'hFF7FFF76;14'd1535:data <=32'hFF66FF85;
14'd1536:data <=32'h0015FFA9;14'd1537:data <=32'hFFFAFF84;14'd1538:data <=32'hFFCAFF77;
14'd1539:data <=32'hFF4BFFD0;14'd1540:data <=32'hFF180007;14'd1541:data <=32'hFF2C002F;
14'd1542:data <=32'hFF47004E;14'd1543:data <=32'hFF670062;14'd1544:data <=32'hFF85006B;
14'd1545:data <=32'hFFA1006E;14'd1546:data <=32'hFFB9006C;14'd1547:data <=32'hFFCE0064;
14'd1548:data <=32'hFFDF0058;14'd1549:data <=32'hFFEB0049;14'd1550:data <=32'hFFED0039;
14'd1551:data <=32'hFFE9002A;14'd1552:data <=32'hFFDD0020;14'd1553:data <=32'hFFCD001F;
14'd1554:data <=32'hFFBD0027;14'd1555:data <=32'hFFB2003A;14'd1556:data <=32'hFFB10051;
14'd1557:data <=32'hFFB9006A;14'd1558:data <=32'hFFCC007E;14'd1559:data <=32'hFFE6008B;
14'd1560:data <=32'h0002008F;14'd1561:data <=32'h001E008A;14'd1562:data <=32'h0036007E;
14'd1563:data <=32'h0047006D;14'd1564:data <=32'h0054005A;14'd1565:data <=32'h005A0046;
14'd1566:data <=32'h005D0032;14'd1567:data <=32'h005B001D;14'd1568:data <=32'h0055000B;
14'd1569:data <=32'h0048FFFC;14'd1570:data <=32'h0038FFF2;14'd1571:data <=32'h0026FFEE;
14'd1572:data <=32'h0013FFF2;14'd1573:data <=32'h0005FFFC;14'd1574:data <=32'hFFFC000C;
14'd1575:data <=32'hFFFA001D;14'd1576:data <=32'h0000002E;14'd1577:data <=32'h000C003A;
14'd1578:data <=32'h00190041;14'd1579:data <=32'h00280043;14'd1580:data <=32'h00350043;
14'd1581:data <=32'h00400041;14'd1582:data <=32'h004A003F;14'd1583:data <=32'h0056003E;
14'd1584:data <=32'h0063003B;14'd1585:data <=32'h00760037;14'd1586:data <=32'h0089002D;
14'd1587:data <=32'h009F001F;14'd1588:data <=32'h00B10006;14'd1589:data <=32'h00BFFFE9;
14'd1590:data <=32'h00C5FFC7;14'd1591:data <=32'h00C5FFA1;14'd1592:data <=32'h00BDFF7C;
14'd1593:data <=32'h00ADFF58;14'd1594:data <=32'h0096FF35;14'd1595:data <=32'h0078FF15;
14'd1596:data <=32'h0051FEFA;14'd1597:data <=32'h0021FEE4;14'd1598:data <=32'hFFEAFED9;
14'd1599:data <=32'hFFB0FEDE;14'd1600:data <=32'h0016FFAE;14'd1601:data <=32'h0010FF8E;
14'd1602:data <=32'hFFF9FF63;14'd1603:data <=32'hFF77FF15;14'd1604:data <=32'hFF1CFF51;
14'd1605:data <=32'hFF0FFF89;14'd1606:data <=32'hFF10FFBD;14'd1607:data <=32'hFF1EFFEA;
14'd1608:data <=32'hFF31000F;14'd1609:data <=32'hFF4A002B;14'd1610:data <=32'hFF650040;
14'd1611:data <=32'hFF81004D;14'd1612:data <=32'hFF9D0051;14'd1613:data <=32'hFFB7004F;
14'd1614:data <=32'hFFCC0045;14'd1615:data <=32'hFFDA0036;14'd1616:data <=32'hFFDD0024;
14'd1617:data <=32'hFFDA0017;14'd1618:data <=32'hFFCF000F;14'd1619:data <=32'hFFC20011;
14'd1620:data <=32'hFFB70019;14'd1621:data <=32'hFFB30027;14'd1622:data <=32'hFFB50035;
14'd1623:data <=32'hFFBC0042;14'd1624:data <=32'hFFC8004B;14'd1625:data <=32'hFFD3004F;
14'd1626:data <=32'hFFDE0050;14'd1627:data <=32'hFFE6004E;14'd1628:data <=32'hFFEB004D;
14'd1629:data <=32'hFFF1004D;14'd1630:data <=32'hFFF7004D;14'd1631:data <=32'hFFFE004E;
14'd1632:data <=32'h0005004D;14'd1633:data <=32'h000C004A;14'd1634:data <=32'h00120045;
14'd1635:data <=32'h00160040;14'd1636:data <=32'h0018003B;14'd1637:data <=32'h00190038;
14'd1638:data <=32'h001A0036;14'd1639:data <=32'h001D0035;14'd1640:data <=32'h00210032;
14'd1641:data <=32'h0024002E;14'd1642:data <=32'h00260028;14'd1643:data <=32'h00230020;
14'd1644:data <=32'h001D001B;14'd1645:data <=32'h00130018;14'd1646:data <=32'h0007001E;
14'd1647:data <=32'hFFFD002B;14'd1648:data <=32'hFFF8003F;14'd1649:data <=32'hFFFD0056;
14'd1650:data <=32'h000D006E;14'd1651:data <=32'h00270082;14'd1652:data <=32'h0049008C;
14'd1653:data <=32'h0070008E;14'd1654:data <=32'h00980082;14'd1655:data <=32'h00BE006C;
14'd1656:data <=32'h00DD004C;14'd1657:data <=32'h00F80025;14'd1658:data <=32'h010AFFF6;
14'd1659:data <=32'h0112FFC1;14'd1660:data <=32'h010EFF88;14'd1661:data <=32'h00FAFF4E;
14'd1662:data <=32'h00D7FF19;14'd1663:data <=32'h00A5FEEC;14'd1664:data <=32'h007AFF6C;
14'd1665:data <=32'h006BFF44;14'd1666:data <=32'h0063FF23;14'd1667:data <=32'h006AFEFA;
14'd1668:data <=32'h0001FF06;14'd1669:data <=32'hFFDDFF16;14'd1670:data <=32'hFFC0FF29;
14'd1671:data <=32'hFFABFF3E;14'd1672:data <=32'hFF98FF53;14'd1673:data <=32'hFF88FF68;
14'd1674:data <=32'hFF7BFF7C;14'd1675:data <=32'hFF70FF93;14'd1676:data <=32'hFF6AFFAB;
14'd1677:data <=32'hFF69FFC2;14'd1678:data <=32'hFF6BFFD7;14'd1679:data <=32'hFF70FFE9;
14'd1680:data <=32'hFF76FFF8;14'd1681:data <=32'hFF7A0004;14'd1682:data <=32'hFF7E0012;
14'd1683:data <=32'hFF840021;14'd1684:data <=32'hFF8C0032;14'd1685:data <=32'hFF9A0041;
14'd1686:data <=32'hFFAD004E;14'd1687:data <=32'hFFC40053;14'd1688:data <=32'hFFDB0051;
14'd1689:data <=32'hFFF00047;14'd1690:data <=32'hFFFD0036;14'd1691:data <=32'h00020023;
14'd1692:data <=32'hFFFE0012;14'd1693:data <=32'hFFF50004;14'd1694:data <=32'hFFE8FFFE;
14'd1695:data <=32'hFFDAFFFD;14'd1696:data <=32'hFFCE0002;14'd1697:data <=32'hFFC4000A;
14'd1698:data <=32'hFFBC0014;14'd1699:data <=32'hFFB90022;14'd1700:data <=32'hFFB80030;
14'd1701:data <=32'hFFBB003F;14'd1702:data <=32'hFFC3004D;14'd1703:data <=32'hFFCD005A;
14'd1704:data <=32'hFFDE0063;14'd1705:data <=32'hFFF00067;14'd1706:data <=32'h00020064;
14'd1707:data <=32'h00110059;14'd1708:data <=32'h0019004C;14'd1709:data <=32'h001A003E;
14'd1710:data <=32'h00130033;14'd1711:data <=32'h0008002E;14'd1712:data <=32'hFFFB0032;
14'd1713:data <=32'hFFF2003E;14'd1714:data <=32'hFFF00050;14'd1715:data <=32'hFFF50064;
14'd1716:data <=32'h00030076;14'd1717:data <=32'h00180086;14'd1718:data <=32'h0032008E;
14'd1719:data <=32'h004D0090;14'd1720:data <=32'h006B008C;14'd1721:data <=32'h00880081;
14'd1722:data <=32'h00A40070;14'd1723:data <=32'h00BF0059;14'd1724:data <=32'h00D3003A;
14'd1725:data <=32'h00E30016;14'd1726:data <=32'h00E9FFEB;14'd1727:data <=32'h00E4FFC1;
14'd1728:data <=32'h0114FFF1;14'd1729:data <=32'h0123FFB0;14'd1730:data <=32'h0116FF82;
14'd1731:data <=32'h00C5FFB9;14'd1732:data <=32'h0080FFB4;14'd1733:data <=32'h007CFFAD;
14'd1734:data <=32'h007CFFA4;14'd1735:data <=32'h007CFF96;14'd1736:data <=32'h007AFF80;
14'd1737:data <=32'h006FFF69;14'd1738:data <=32'h005DFF50;14'd1739:data <=32'h0042FF3B;
14'd1740:data <=32'h0022FF2D;14'd1741:data <=32'hFFFFFF27;14'd1742:data <=32'hFFDBFF29;
14'd1743:data <=32'hFFB7FF31;14'd1744:data <=32'hFF95FF40;14'd1745:data <=32'hFF76FF57;
14'd1746:data <=32'hFF59FF73;14'd1747:data <=32'hFF44FF98;14'd1748:data <=32'hFF38FFC3;
14'd1749:data <=32'hFF38FFEF;14'd1750:data <=32'hFF46001B;14'd1751:data <=32'hFF61003F;
14'd1752:data <=32'hFF830059;14'd1753:data <=32'hFFAB0064;14'd1754:data <=32'hFFD10063;
14'd1755:data <=32'hFFF10055;14'd1756:data <=32'h00060041;14'd1757:data <=32'h00130028;
14'd1758:data <=32'h00170010;14'd1759:data <=32'h0013FFFB;14'd1760:data <=32'h000AFFE9;
14'd1761:data <=32'hFFFDFFDC;14'd1762:data <=32'hFFEEFFD3;14'd1763:data <=32'hFFDDFFCE;
14'd1764:data <=32'hFFC9FFCE;14'd1765:data <=32'hFFB7FFD4;14'd1766:data <=32'hFFA6FFDF;
14'd1767:data <=32'hFF99FFF0;14'd1768:data <=32'hFF910003;14'd1769:data <=32'hFF8F0018;
14'd1770:data <=32'hFF91002A;14'd1771:data <=32'hFF980039;14'd1772:data <=32'hFFA10044;
14'd1773:data <=32'hFFA8004D;14'd1774:data <=32'hFFAD0055;14'd1775:data <=32'hFFB0005E;
14'd1776:data <=32'hFFB3006B;14'd1777:data <=32'hFFBB007B;14'd1778:data <=32'hFFC7008C;
14'd1779:data <=32'hFFD9009C;14'd1780:data <=32'hFFF100A8;14'd1781:data <=32'h000D00AE;
14'd1782:data <=32'h002B00AC;14'd1783:data <=32'h004600A2;14'd1784:data <=32'h005D0094;
14'd1785:data <=32'h006F0081;14'd1786:data <=32'h007D006D;14'd1787:data <=32'h0086005A;
14'd1788:data <=32'h008D0046;14'd1789:data <=32'h00900032;14'd1790:data <=32'h008E001E;
14'd1791:data <=32'h0089000B;14'd1792:data <=32'h00BB00B5;14'd1793:data <=32'h00F30093;
14'd1794:data <=32'h0108005A;14'd1795:data <=32'h007F0006;14'd1796:data <=32'h003F0014;
14'd1797:data <=32'h00460023;14'd1798:data <=32'h0058002E;14'd1799:data <=32'h00700031;
14'd1800:data <=32'h008D0027;14'd1801:data <=32'h00A60010;14'd1802:data <=32'h00B6FFF1;
14'd1803:data <=32'h00BDFFCD;14'd1804:data <=32'h00B9FFA5;14'd1805:data <=32'h00ACFF80;
14'd1806:data <=32'h0096FF60;14'd1807:data <=32'h0079FF44;14'd1808:data <=32'h0056FF2F;
14'd1809:data <=32'h002EFF20;14'd1810:data <=32'h0001FF1C;14'd1811:data <=32'hFFD5FF23;
14'd1812:data <=32'hFFAAFF36;14'd1813:data <=32'hFF86FF54;14'd1814:data <=32'hFF6EFF7B;
14'd1815:data <=32'hFF62FFA6;14'd1816:data <=32'hFF65FFCE;14'd1817:data <=32'hFF72FFF1;
14'd1818:data <=32'hFF85000B;14'd1819:data <=32'hFF9D001B;14'd1820:data <=32'hFFB30024;
14'd1821:data <=32'hFFC80026;14'd1822:data <=32'hFFD90024;14'd1823:data <=32'hFFE70021;
14'd1824:data <=32'hFFF5001B;14'd1825:data <=32'h00000012;14'd1826:data <=32'h000B0007;
14'd1827:data <=32'h0012FFF8;14'd1828:data <=32'h0014FFE7;14'd1829:data <=32'h0011FFD5;
14'd1830:data <=32'h0008FFC3;14'd1831:data <=32'hFFF9FFB5;14'd1832:data <=32'hFFE7FFAB;
14'd1833:data <=32'hFFD3FFA5;14'd1834:data <=32'hFFBDFFA4;14'd1835:data <=32'hFFA7FFA6;
14'd1836:data <=32'hFF90FFAD;14'd1837:data <=32'hFF78FFB8;14'd1838:data <=32'hFF60FFCA;
14'd1839:data <=32'hFF48FFE3;14'd1840:data <=32'hFF360003;14'd1841:data <=32'hFF2A002C;
14'd1842:data <=32'hFF2A005A;14'd1843:data <=32'hFF38008A;14'd1844:data <=32'hFF5200B6;
14'd1845:data <=32'hFF7A00D9;14'd1846:data <=32'hFFA900EF;14'd1847:data <=32'hFFDA00F8;
14'd1848:data <=32'h000C00F2;14'd1849:data <=32'h003600E4;14'd1850:data <=32'h005900CD;
14'd1851:data <=32'h007400B0;14'd1852:data <=32'h00860090;14'd1853:data <=32'h00910071;
14'd1854:data <=32'h00930050;14'd1855:data <=32'h008E0032;14'd1856:data <=32'h002A00A2;
14'd1857:data <=32'h004D00A7;14'd1858:data <=32'h00790096;14'd1859:data <=32'h0095002D;
14'd1860:data <=32'h004C002B;14'd1861:data <=32'h00470032;14'd1862:data <=32'h004A003B;
14'd1863:data <=32'h00550043;14'd1864:data <=32'h00660045;14'd1865:data <=32'h007B003E;
14'd1866:data <=32'h008B002D;14'd1867:data <=32'h00980018;14'd1868:data <=32'h009D0000;
14'd1869:data <=32'h009DFFE9;14'd1870:data <=32'h0098FFD3;14'd1871:data <=32'h0090FFBE;
14'd1872:data <=32'h0085FFAB;14'd1873:data <=32'h0077FF99;14'd1874:data <=32'h0065FF88;
14'd1875:data <=32'h004FFF7D;14'd1876:data <=32'h0037FF76;14'd1877:data <=32'h001DFF76;
14'd1878:data <=32'h0007FF7D;14'd1879:data <=32'hFFF5FF8A;14'd1880:data <=32'hFFEAFF97;
14'd1881:data <=32'hFFE4FFA4;14'd1882:data <=32'hFFE2FFAC;14'd1883:data <=32'hFFE0FFB3;
14'd1884:data <=32'hFFDDFFB7;14'd1885:data <=32'hFFD6FFBB;14'd1886:data <=32'hFFCEFFC2;
14'd1887:data <=32'hFFC7FFCD;14'd1888:data <=32'hFFC3FFDA;14'd1889:data <=32'hFFC5FFEB;
14'd1890:data <=32'hFFCDFFFA;14'd1891:data <=32'hFFDA0005;14'd1892:data <=32'hFFEB000B;
14'd1893:data <=32'hFFFD0009;14'd1894:data <=32'h000F0001;14'd1895:data <=32'h001CFFF5;
14'd1896:data <=32'h0025FFE2;14'd1897:data <=32'h0028FFCD;14'd1898:data <=32'h0027FFB7;
14'd1899:data <=32'h001EFF9F;14'd1900:data <=32'h000EFF87;14'd1901:data <=32'hFFF5FF72;
14'd1902:data <=32'hFFD5FF63;14'd1903:data <=32'hFFADFF5C;14'd1904:data <=32'hFF80FF61;
14'd1905:data <=32'hFF53FF73;14'd1906:data <=32'hFF2DFF95;14'd1907:data <=32'hFF0FFFC2;
14'd1908:data <=32'hFF01FFF6;14'd1909:data <=32'hFF00002C;14'd1910:data <=32'hFF0F005D;
14'd1911:data <=32'hFF280087;14'd1912:data <=32'hFF4900A8;14'd1913:data <=32'hFF6C00BF;
14'd1914:data <=32'hFF9200CD;14'd1915:data <=32'hFFB500D4;14'd1916:data <=32'hFFD800D5;
14'd1917:data <=32'hFFF800D1;14'd1918:data <=32'h001500C6;14'd1919:data <=32'h002E00B6;
14'd1920:data <=32'h00250088;14'd1921:data <=32'h00320085;14'd1922:data <=32'h003F008C;
14'd1923:data <=32'h004B00C6;14'd1924:data <=32'h002300BD;14'd1925:data <=32'h003900BC;
14'd1926:data <=32'h005300B8;14'd1927:data <=32'h006F00AF;14'd1928:data <=32'h008E009E;
14'd1929:data <=32'h00A80083;14'd1930:data <=32'h00BC0061;14'd1931:data <=32'h00C4003A;
14'd1932:data <=32'h00C20013;14'd1933:data <=32'h00B4FFF2;14'd1934:data <=32'h00A0FFD7;
14'd1935:data <=32'h008AFFC4;14'd1936:data <=32'h0072FFB9;14'd1937:data <=32'h005DFFB4;
14'd1938:data <=32'h0049FFB3;14'd1939:data <=32'h0037FFB7;14'd1940:data <=32'h0027FFBD;
14'd1941:data <=32'h001BFFC7;14'd1942:data <=32'h0015FFD4;14'd1943:data <=32'h0014FFE1;
14'd1944:data <=32'h001AFFED;14'd1945:data <=32'h0026FFF3;14'd1946:data <=32'h0033FFF2;
14'd1947:data <=32'h003FFFEA;14'd1948:data <=32'h0046FFDA;14'd1949:data <=32'h0046FFC8;
14'd1950:data <=32'h003CFFB7;14'd1951:data <=32'h002DFFAB;14'd1952:data <=32'h001BFFA6;
14'd1953:data <=32'h0008FFA9;14'd1954:data <=32'hFFFAFFB1;14'd1955:data <=32'hFFF1FFBD;
14'd1956:data <=32'hFFEDFFCA;14'd1957:data <=32'hFFEFFFD6;14'd1958:data <=32'hFFF4FFDD;
14'd1959:data <=32'hFFFCFFE3;14'd1960:data <=32'h0005FFE4;14'd1961:data <=32'h000EFFE3;
14'd1962:data <=32'h0018FFDD;14'd1963:data <=32'h0020FFD3;14'd1964:data <=32'h0026FFC5;
14'd1965:data <=32'h0028FFB2;14'd1966:data <=32'h0023FF9D;14'd1967:data <=32'h0015FF88;
14'd1968:data <=32'hFFFFFF76;14'd1969:data <=32'hFFE3FF6B;14'd1970:data <=32'hFFC4FF69;
14'd1971:data <=32'hFFA5FF70;14'd1972:data <=32'hFF8AFF7F;14'd1973:data <=32'hFF75FF93;
14'd1974:data <=32'hFF67FFA9;14'd1975:data <=32'hFF5EFFBE;14'd1976:data <=32'hFF57FFD2;
14'd1977:data <=32'hFF51FFE2;14'd1978:data <=32'hFF4BFFF5;14'd1979:data <=32'hFF450009;
14'd1980:data <=32'hFF400020;14'd1981:data <=32'hFF3E003A;14'd1982:data <=32'hFF420057;
14'd1983:data <=32'hFF4B0074;14'd1984:data <=32'hFFC800B1;14'd1985:data <=32'hFFDD00B2;
14'd1986:data <=32'hFFDD00A8;14'd1987:data <=32'hFF6100A7;14'd1988:data <=32'hFF3B00C9;
14'd1989:data <=32'hFF5D00F1;14'd1990:data <=32'hFF8A0113;14'd1991:data <=32'hFFC0012A;
14'd1992:data <=32'hFFFF0133;14'd1993:data <=32'h003F012A;14'd1994:data <=32'h007A010F;
14'd1995:data <=32'h00AA00E5;14'd1996:data <=32'h00CB00B2;14'd1997:data <=32'h00DC007B;
14'd1998:data <=32'h00DC0047;14'd1999:data <=32'h00D10018;14'd2000:data <=32'h00BCFFF2;
14'd2001:data <=32'h00A3FFD5;14'd2002:data <=32'h0086FFC0;14'd2003:data <=32'h0067FFB5;
14'd2004:data <=32'h0048FFB0;14'd2005:data <=32'h002CFFB5;14'd2006:data <=32'h0012FFC3;
14'd2007:data <=32'h0002FFD6;14'd2008:data <=32'hFFFAFFEC;14'd2009:data <=32'hFFFC0002;
14'd2010:data <=32'h00070014;14'd2011:data <=32'h0017001E;14'd2012:data <=32'h00290020;
14'd2013:data <=32'h0038001B;14'd2014:data <=32'h00430011;14'd2015:data <=32'h00480004;
14'd2016:data <=32'h0049FFFA;14'd2017:data <=32'h0047FFF2;14'd2018:data <=32'h0045FFED;
14'd2019:data <=32'h0045FFE9;14'd2020:data <=32'h0045FFE4;14'd2021:data <=32'h0047FFDF;
14'd2022:data <=32'h0049FFD7;14'd2023:data <=32'h0049FFCD;14'd2024:data <=32'h0045FFC3;
14'd2025:data <=32'h003FFFB8;14'd2026:data <=32'h0038FFB1;14'd2027:data <=32'h0030FFAA;
14'd2028:data <=32'h0028FFA6;14'd2029:data <=32'h001FFFA2;14'd2030:data <=32'h0017FF9E;
14'd2031:data <=32'h000DFF99;14'd2032:data <=32'h0002FF97;14'd2033:data <=32'hFFF5FF97;
14'd2034:data <=32'hFFE9FF9A;14'd2035:data <=32'hFFDDFFA2;14'd2036:data <=32'hFFD7FFAB;
14'd2037:data <=32'hFFD7FFB4;14'd2038:data <=32'hFFDCFFBA;14'd2039:data <=32'hFFE3FFB7;
14'd2040:data <=32'hFFE8FFAF;14'd2041:data <=32'hFFE7FFA0;14'd2042:data <=32'hFFDDFF8E;
14'd2043:data <=32'hFFC8FF7E;14'd2044:data <=32'hFFADFF74;14'd2045:data <=32'hFF89FF72;
14'd2046:data <=32'hFF65FF7B;14'd2047:data <=32'hFF42FF8F;14'd2048:data <=32'hFF50001B;
14'd2049:data <=32'hFF4B002E;14'd2050:data <=32'hFF53002D;14'd2051:data <=32'hFF39FFCB;
14'd2052:data <=32'hFEEAFFF1;14'd2053:data <=32'hFEE10029;14'd2054:data <=32'hFEE80063;
14'd2055:data <=32'hFEFD009C;14'd2056:data <=32'hFF2300CF;14'd2057:data <=32'hFF5600F5;
14'd2058:data <=32'hFF8F010B;14'd2059:data <=32'hFFCA010F;14'd2060:data <=32'h00000105;
14'd2061:data <=32'h002C00EF;14'd2062:data <=32'h004F00D3;14'd2063:data <=32'h006800B4;
14'd2064:data <=32'h00790095;14'd2065:data <=32'h00830078;14'd2066:data <=32'h0087005A;
14'd2067:data <=32'h0087003E;14'd2068:data <=32'h00810024;14'd2069:data <=32'h0075000D;
14'd2070:data <=32'h0066FFFC;14'd2071:data <=32'h0054FFF1;14'd2072:data <=32'h0042FFEC;
14'd2073:data <=32'h0032FFED;14'd2074:data <=32'h0028FFF1;14'd2075:data <=32'h0020FFF7;
14'd2076:data <=32'h001BFFFB;14'd2077:data <=32'h0017FFFE;14'd2078:data <=32'h00120000;
14'd2079:data <=32'h000C0005;14'd2080:data <=32'h0007000E;14'd2081:data <=32'h0004001A;
14'd2082:data <=32'h00070029;14'd2083:data <=32'h00100039;14'd2084:data <=32'h00210045;
14'd2085:data <=32'h0037004A;14'd2086:data <=32'h00510049;14'd2087:data <=32'h0069003E;
14'd2088:data <=32'h007E002C;14'd2089:data <=32'h008D0014;14'd2090:data <=32'h0094FFF8;
14'd2091:data <=32'h0095FFDD;14'd2092:data <=32'h008FFFC3;14'd2093:data <=32'h0084FFAB;
14'd2094:data <=32'h0074FF95;14'd2095:data <=32'h005FFF84;14'd2096:data <=32'h0047FF78;
14'd2097:data <=32'h002CFF72;14'd2098:data <=32'h0012FF74;14'd2099:data <=32'hFFFBFF7F;
14'd2100:data <=32'hFFEAFF90;14'd2101:data <=32'hFFE1FFA4;14'd2102:data <=32'hFFE3FFB8;
14'd2103:data <=32'hFFEEFFC4;14'd2104:data <=32'hFFFCFFC8;14'd2105:data <=32'h000DFFC1;
14'd2106:data <=32'h0017FFB1;14'd2107:data <=32'h0019FF9C;14'd2108:data <=32'h0010FF84;
14'd2109:data <=32'hFFFEFF6E;14'd2110:data <=32'hFFE4FF5F;14'd2111:data <=32'hFFC4FF56;
14'd2112:data <=32'hFFCFFF71;14'd2113:data <=32'hFFADFF61;14'd2114:data <=32'hFF98FF64;
14'd2115:data <=32'hFFABFF89;14'd2116:data <=32'hFF58FF90;14'd2117:data <=32'hFF44FFAA;
14'd2118:data <=32'hFF36FFCA;14'd2119:data <=32'hFF2FFFEE;14'd2120:data <=32'hFF320012;
14'd2121:data <=32'hFF3F0034;14'd2122:data <=32'hFF53004E;14'd2123:data <=32'hFF6A0060;
14'd2124:data <=32'hFF80006A;14'd2125:data <=32'hFF93006E;14'd2126:data <=32'hFFA00071;
14'd2127:data <=32'hFFAB0075;14'd2128:data <=32'hFFB5007B;14'd2129:data <=32'hFFC10084;
14'd2130:data <=32'hFFD0008C;14'd2131:data <=32'hFFE30092;14'd2132:data <=32'hFFF90093;
14'd2133:data <=32'h0010008F;14'd2134:data <=32'h00230086;14'd2135:data <=32'h0035007B;
14'd2136:data <=32'h0043006D;14'd2137:data <=32'h004E005D;14'd2138:data <=32'h0057004B;
14'd2139:data <=32'h005E0037;14'd2140:data <=32'h005E0021;14'd2141:data <=32'h0059000A;
14'd2142:data <=32'h004CFFF5;14'd2143:data <=32'h0038FFE5;14'd2144:data <=32'h001EFFDD;
14'd2145:data <=32'h0003FFE0;14'd2146:data <=32'hFFEBFFED;14'd2147:data <=32'hFFDA0004;
14'd2148:data <=32'hFFD3001F;14'd2149:data <=32'hFFD6003D;14'd2150:data <=32'hFFE50057;
14'd2151:data <=32'hFFFC006A;14'd2152:data <=32'h00170075;14'd2153:data <=32'h00340078;
14'd2154:data <=32'h00500073;14'd2155:data <=32'h00690067;14'd2156:data <=32'h007F0057;
14'd2157:data <=32'h00910042;14'd2158:data <=32'h009F0029;14'd2159:data <=32'h00A6000F;
14'd2160:data <=32'h00A9FFF2;14'd2161:data <=32'h00A3FFD7;14'd2162:data <=32'h0098FFBE;
14'd2163:data <=32'h0087FFAB;14'd2164:data <=32'h0075FF9F;14'd2165:data <=32'h0065FF98;
14'd2166:data <=32'h0058FF97;14'd2167:data <=32'h0050FF95;14'd2168:data <=32'h004CFF91;
14'd2169:data <=32'h004AFF89;14'd2170:data <=32'h0044FF7C;14'd2171:data <=32'h003AFF6B;
14'd2172:data <=32'h0028FF5B;14'd2173:data <=32'h0011FF4F;14'd2174:data <=32'hFFF6FF4A;
14'd2175:data <=32'hFFD9FF4B;14'd2176:data <=32'h0063FFB0;14'd2177:data <=32'h0061FF7E;
14'd2178:data <=32'h0042FF57;14'd2179:data <=32'hFFB5FF78;14'd2180:data <=32'hFF6BFF85;
14'd2181:data <=32'hFF64FFA4;14'd2182:data <=32'hFF62FFC1;14'd2183:data <=32'hFF67FFDD;
14'd2184:data <=32'hFF73FFF6;14'd2185:data <=32'hFF840009;14'd2186:data <=32'hFF9A0013;
14'd2187:data <=32'hFFAF0014;14'd2188:data <=32'hFFBE000C;14'd2189:data <=32'hFFC5FFFE;
14'd2190:data <=32'hFFC2FFF0;14'd2191:data <=32'hFFB4FFE7;14'd2192:data <=32'hFFA3FFE6;
14'd2193:data <=32'hFF90FFEF;14'd2194:data <=32'hFF800000;14'd2195:data <=32'hFF790017;
14'd2196:data <=32'hFF780032;14'd2197:data <=32'hFF7F004B;14'd2198:data <=32'hFF8C0061;
14'd2199:data <=32'hFF9E0074;14'd2200:data <=32'hFFB20083;14'd2201:data <=32'hFFCC008D;
14'd2202:data <=32'hFFE70091;14'd2203:data <=32'h0004008F;14'd2204:data <=32'h00200083;
14'd2205:data <=32'h00380071;14'd2206:data <=32'h00460056;14'd2207:data <=32'h004C003A;
14'd2208:data <=32'h0048001E;14'd2209:data <=32'h003A0007;14'd2210:data <=32'h0027FFF9;
14'd2211:data <=32'h0010FFF4;14'd2212:data <=32'hFFFBFFF8;14'd2213:data <=32'hFFEB0003;
14'd2214:data <=32'hFFE10012;14'd2215:data <=32'hFFDD0020;14'd2216:data <=32'hFFDD002F;
14'd2217:data <=32'hFFE0003C;14'd2218:data <=32'hFFE50049;14'd2219:data <=32'hFFEB0056;
14'd2220:data <=32'hFFF50062;14'd2221:data <=32'h0000006E;14'd2222:data <=32'h00120079;
14'd2223:data <=32'h00250080;14'd2224:data <=32'h003C0083;14'd2225:data <=32'h00550082;
14'd2226:data <=32'h006D007B;14'd2227:data <=32'h00840070;14'd2228:data <=32'h00990062;
14'd2229:data <=32'h00AE0051;14'd2230:data <=32'h00C2003D;14'd2231:data <=32'h00D50024;
14'd2232:data <=32'h00E60003;14'd2233:data <=32'h00F3FFDB;14'd2234:data <=32'h00F5FFAD;
14'd2235:data <=32'h00ECFF7B;14'd2236:data <=32'h00D4FF4B;14'd2237:data <=32'h00AEFF20;
14'd2238:data <=32'h007EFF02;14'd2239:data <=32'h0048FEF2;14'd2240:data <=32'h0058FFE5;
14'd2241:data <=32'h0070FFC6;14'd2242:data <=32'h0079FF8F;14'd2243:data <=32'h0016FF0D;
14'd2244:data <=32'hFFB2FF13;14'd2245:data <=32'hFF8FFF33;14'd2246:data <=32'hFF77FF59;
14'd2247:data <=32'hFF69FF81;14'd2248:data <=32'hFF66FFA9;14'd2249:data <=32'hFF6FFFCE;
14'd2250:data <=32'hFF83FFEA;14'd2251:data <=32'hFF9AFFFC;14'd2252:data <=32'hFFB40002;
14'd2253:data <=32'hFFCAFFFC;14'd2254:data <=32'hFFD7FFEF;14'd2255:data <=32'hFFD9FFE0;
14'd2256:data <=32'hFFD2FFD3;14'd2257:data <=32'hFFC6FFCC;14'd2258:data <=32'hFFB7FFCD;
14'd2259:data <=32'hFFA9FFD2;14'd2260:data <=32'hFF9EFFDE;14'd2261:data <=32'hFF97FFEB;
14'd2262:data <=32'hFF93FFF9;14'd2263:data <=32'hFF920007;14'd2264:data <=32'hFF920016;
14'd2265:data <=32'hFF960025;14'd2266:data <=32'hFF9C0034;14'd2267:data <=32'hFFA60042;
14'd2268:data <=32'hFFB5004D;14'd2269:data <=32'hFFC60052;14'd2270:data <=32'hFFD60052;
14'd2271:data <=32'hFFE4004E;14'd2272:data <=32'hFFEF0046;14'd2273:data <=32'hFFF4003D;
14'd2274:data <=32'hFFF60036;14'd2275:data <=32'hFFF50032;14'd2276:data <=32'hFFF50031;
14'd2277:data <=32'hFFF60031;14'd2278:data <=32'hFFF90031;14'd2279:data <=32'hFFFE002E;
14'd2280:data <=32'h00020029;14'd2281:data <=32'h00020020;14'd2282:data <=32'hFFFD0018;
14'd2283:data <=32'hFFF30011;14'd2284:data <=32'hFFE50010;14'd2285:data <=32'hFFD40015;
14'd2286:data <=32'hFFC60023;14'd2287:data <=32'hFFBC0036;14'd2288:data <=32'hFFB7004E;
14'd2289:data <=32'hFFBB006A;14'd2290:data <=32'hFFC60085;14'd2291:data <=32'hFFD7009F;
14'd2292:data <=32'hFFF100B6;14'd2293:data <=32'h001100CA;14'd2294:data <=32'h003900D7;
14'd2295:data <=32'h006800DC;14'd2296:data <=32'h009D00D5;14'd2297:data <=32'h00D100BE;
14'd2298:data <=32'h01020097;14'd2299:data <=32'h01280061;14'd2300:data <=32'h013D0021;
14'd2301:data <=32'h0140FFDE;14'd2302:data <=32'h0131FF9C;14'd2303:data <=32'h0111FF64;
14'd2304:data <=32'h00A0FFD7;14'd2305:data <=32'h00AEFFBA;14'd2306:data <=32'h00C5FF9D;
14'd2307:data <=32'h00EBFF63;14'd2308:data <=32'h008FFF3B;14'd2309:data <=32'h0069FF31;
14'd2310:data <=32'h0044FF2F;14'd2311:data <=32'h0023FF31;14'd2312:data <=32'h0003FF3C;
14'd2313:data <=32'hFFE9FF4C;14'd2314:data <=32'hFFD8FF5F;14'd2315:data <=32'hFFCDFF72;
14'd2316:data <=32'hFFC8FF81;14'd2317:data <=32'hFFC3FF8A;14'd2318:data <=32'hFFBFFF90;
14'd2319:data <=32'hFFB6FF95;14'd2320:data <=32'hFFABFF9D;14'd2321:data <=32'hFF9EFFA8;
14'd2322:data <=32'hFF94FFBA;14'd2323:data <=32'hFF8FFFCE;14'd2324:data <=32'hFF90FFE5;
14'd2325:data <=32'hFF99FFF7;14'd2326:data <=32'hFFA60005;14'd2327:data <=32'hFFB4000C;
14'd2328:data <=32'hFFC1000F;14'd2329:data <=32'hFFCB000E;14'd2330:data <=32'hFFD3000A;
14'd2331:data <=32'hFFD80006;14'd2332:data <=32'hFFDB0001;14'd2333:data <=32'hFFDCFFFC;
14'd2334:data <=32'hFFDBFFF6;14'd2335:data <=32'hFFD7FFF0;14'd2336:data <=32'hFFD0FFEC;
14'd2337:data <=32'hFFC6FFEB;14'd2338:data <=32'hFFB8FFEE;14'd2339:data <=32'hFFADFFF8;
14'd2340:data <=32'hFFA50008;14'd2341:data <=32'hFFA3001A;14'd2342:data <=32'hFFA9002C;
14'd2343:data <=32'hFFB6003A;14'd2344:data <=32'hFFC70042;14'd2345:data <=32'hFFD70043;
14'd2346:data <=32'hFFE5003C;14'd2347:data <=32'hFFED002F;14'd2348:data <=32'hFFEE0022;
14'd2349:data <=32'hFFE80018;14'd2350:data <=32'hFFDC0012;14'd2351:data <=32'hFFCD0012;
14'd2352:data <=32'hFFBF0019;14'd2353:data <=32'hFFB30025;14'd2354:data <=32'hFFA80037;
14'd2355:data <=32'hFFA3004C;14'd2356:data <=32'hFFA20065;14'd2357:data <=32'hFFA80080;
14'd2358:data <=32'hFFB6009F;14'd2359:data <=32'hFFCD00BA;14'd2360:data <=32'hFFEE00D2;
14'd2361:data <=32'h001900E1;14'd2362:data <=32'h004800E4;14'd2363:data <=32'h007800D9;
14'd2364:data <=32'h00A300C1;14'd2365:data <=32'h00C6009D;14'd2366:data <=32'h00DC0075;
14'd2367:data <=32'h00E6004D;14'd2368:data <=32'h00E80078;14'd2369:data <=32'h010F0050;
14'd2370:data <=32'h011F0032;14'd2371:data <=32'h00DE004E;14'd2372:data <=32'h00AE0027;
14'd2373:data <=32'h00B60014;14'd2374:data <=32'h00BDFFFE;14'd2375:data <=32'h00C1FFE5;
14'd2376:data <=32'h00BFFFCB;14'd2377:data <=32'h00BAFFB0;14'd2378:data <=32'h00B1FF97;
14'd2379:data <=32'h00A4FF7E;14'd2380:data <=32'h0094FF65;14'd2381:data <=32'h007EFF4C;
14'd2382:data <=32'h0061FF35;14'd2383:data <=32'h003BFF23;14'd2384:data <=32'h0010FF1B;
14'd2385:data <=32'hFFE1FF1E;14'd2386:data <=32'hFFB5FF31;14'd2387:data <=32'hFF8FFF4E;
14'd2388:data <=32'hFF75FF76;14'd2389:data <=32'hFF6AFFA1;14'd2390:data <=32'hFF6BFFCA;
14'd2391:data <=32'hFF77FFED;14'd2392:data <=32'hFF8B0008;14'd2393:data <=32'hFFA3001B;
14'd2394:data <=32'hFFBB0025;14'd2395:data <=32'hFFD40028;14'd2396:data <=32'hFFEA0025;
14'd2397:data <=32'hFFFE001C;14'd2398:data <=32'h000E000B;14'd2399:data <=32'h0018FFF8;
14'd2400:data <=32'h001AFFE2;14'd2401:data <=32'h0013FFCD;14'd2402:data <=32'h0005FFBB;
14'd2403:data <=32'hFFF1FFAF;14'd2404:data <=32'hFFDAFFAC;14'd2405:data <=32'hFFC4FFB0;
14'd2406:data <=32'hFFB2FFBC;14'd2407:data <=32'hFFA7FFCB;14'd2408:data <=32'hFFA2FFDA;
14'd2409:data <=32'hFFA0FFE6;14'd2410:data <=32'hFFA1FFEF;14'd2411:data <=32'hFFA1FFF6;
14'd2412:data <=32'hFF9EFFFA;14'd2413:data <=32'hFF9A0000;14'd2414:data <=32'hFF930008;
14'd2415:data <=32'hFF8E0014;14'd2416:data <=32'hFF890023;14'd2417:data <=32'hFF890034;
14'd2418:data <=32'hFF8B0045;14'd2419:data <=32'hFF930055;14'd2420:data <=32'hFF9B0064;
14'd2421:data <=32'hFFA60073;14'd2422:data <=32'hFFB20081;14'd2423:data <=32'hFFC0008D;
14'd2424:data <=32'hFFD30098;14'd2425:data <=32'hFFE900A0;14'd2426:data <=32'h000100A3;
14'd2427:data <=32'h001B009F;14'd2428:data <=32'h00300093;14'd2429:data <=32'h00410084;
14'd2430:data <=32'h00480072;14'd2431:data <=32'h004A0066;14'd2432:data <=32'h00420102;
14'd2433:data <=32'h007C0103;14'd2434:data <=32'h00A500E5;14'd2435:data <=32'h0046007A;
14'd2436:data <=32'h00170071;14'd2437:data <=32'h00280081;14'd2438:data <=32'h0040008B;
14'd2439:data <=32'h005E008E;14'd2440:data <=32'h007E0089;14'd2441:data <=32'h009C007C;
14'd2442:data <=32'h00BA0067;14'd2443:data <=32'h00D3004A;14'd2444:data <=32'h00E90026;
14'd2445:data <=32'h00F6FFF9;14'd2446:data <=32'h00F7FFC8;14'd2447:data <=32'h00EBFF96;
14'd2448:data <=32'h00CFFF65;14'd2449:data <=32'h00A7FF40;14'd2450:data <=32'h0075FF27;
14'd2451:data <=32'h0040FF1F;14'd2452:data <=32'h000EFF25;14'd2453:data <=32'hFFE4FF39;
14'd2454:data <=32'hFFC3FF55;14'd2455:data <=32'hFFAEFF74;14'd2456:data <=32'hFFA2FF93;
14'd2457:data <=32'hFF9DFFB1;14'd2458:data <=32'hFF9FFFCC;14'd2459:data <=32'hFFA6FFE4;
14'd2460:data <=32'hFFB2FFFA;14'd2461:data <=32'hFFC3000A;14'd2462:data <=32'hFFD70015;
14'd2463:data <=32'hFFED001A;14'd2464:data <=32'h00010017;14'd2465:data <=32'h0013000C;
14'd2466:data <=32'h0020FFFE;14'd2467:data <=32'h0028FFEC;14'd2468:data <=32'h0029FFDB;
14'd2469:data <=32'h0026FFCC;14'd2470:data <=32'h0021FFBF;14'd2471:data <=32'h001AFFB2;
14'd2472:data <=32'h0013FFA6;14'd2473:data <=32'h0009FF99;14'd2474:data <=32'hFFFCFF8B;
14'd2475:data <=32'hFFE8FF7D;14'd2476:data <=32'hFFCFFF73;14'd2477:data <=32'hFFB0FF70;
14'd2478:data <=32'hFF8DFF75;14'd2479:data <=32'hFF6AFF85;14'd2480:data <=32'hFF4AFF9F;
14'd2481:data <=32'hFF34FFC1;14'd2482:data <=32'hFF26FFE9;14'd2483:data <=32'hFF240013;
14'd2484:data <=32'hFF2A003B;14'd2485:data <=32'hFF39005F;14'd2486:data <=32'hFF4F007E;
14'd2487:data <=32'hFF6A0099;14'd2488:data <=32'hFF8B00AD;14'd2489:data <=32'hFFAE00B8;
14'd2490:data <=32'hFFD400BA;14'd2491:data <=32'hFFF800B3;14'd2492:data <=32'h001500A1;
14'd2493:data <=32'h002B0088;14'd2494:data <=32'h0034006C;14'd2495:data <=32'h00310052;
14'd2496:data <=32'hFFB0009B;14'd2497:data <=32'hFFC300B8;14'd2498:data <=32'hFFED00C6;
14'd2499:data <=32'h002B006C;14'd2500:data <=32'hFFF0005C;14'd2501:data <=32'hFFF2006B;
14'd2502:data <=32'hFFFA007A;14'd2503:data <=32'h000A0087;14'd2504:data <=32'h001C008F;
14'd2505:data <=32'h00330092;14'd2506:data <=32'h004A0092;14'd2507:data <=32'h0064008D;
14'd2508:data <=32'h007E0083;14'd2509:data <=32'h00980070;14'd2510:data <=32'h00AE0055;
14'd2511:data <=32'h00BD0035;14'd2512:data <=32'h00C30010;14'd2513:data <=32'h00BEFFEB;
14'd2514:data <=32'h00ADFFCB;14'd2515:data <=32'h0098FFB2;14'd2516:data <=32'h007FFFA2;
14'd2517:data <=32'h0066FF9C;14'd2518:data <=32'h0052FF9A;14'd2519:data <=32'h0041FF9A;
14'd2520:data <=32'h0035FF9B;14'd2521:data <=32'h0027FF9B;14'd2522:data <=32'h001AFF9C;
14'd2523:data <=32'h000CFF9F;14'd2524:data <=32'hFFFDFFA5;14'd2525:data <=32'hFFF0FFAF;
14'd2526:data <=32'hFFE6FFBC;14'd2527:data <=32'hFFE1FFCA;14'd2528:data <=32'hFFE0FFD9;
14'd2529:data <=32'hFFE3FFE7;14'd2530:data <=32'hFFEAFFF2;14'd2531:data <=32'hFFF2FFFC;
14'd2532:data <=32'hFFFE0004;14'd2533:data <=32'h000B0008;14'd2534:data <=32'h001A000B;
14'd2535:data <=32'h002C0007;14'd2536:data <=32'h0041FFFE;14'd2537:data <=32'h0053FFEC;
14'd2538:data <=32'h0061FFD2;14'd2539:data <=32'h0067FFB0;14'd2540:data <=32'h0062FF8A;
14'd2541:data <=32'h004FFF65;14'd2542:data <=32'h0030FF44;14'd2543:data <=32'h0006FF2F;
14'd2544:data <=32'hFFD6FF26;14'd2545:data <=32'hFFA5FF2B;14'd2546:data <=32'hFF78FF3C;
14'd2547:data <=32'hFF52FF57;14'd2548:data <=32'hFF34FF7B;14'd2549:data <=32'hFF1FFFA2;
14'd2550:data <=32'hFF13FFCC;14'd2551:data <=32'hFF0FFFF7;14'd2552:data <=32'hFF160021;
14'd2553:data <=32'hFF260049;14'd2554:data <=32'hFF3D006B;14'd2555:data <=32'hFF5C0084;
14'd2556:data <=32'hFF7E0092;14'd2557:data <=32'hFF9F0096;14'd2558:data <=32'hFFBA0090;
14'd2559:data <=32'hFFCD0085;14'd2560:data <=32'hFFCD0053;14'd2561:data <=32'hFFC70056;
14'd2562:data <=32'hFFC5006C;14'd2563:data <=32'hFFC600AE;14'd2564:data <=32'hFFA100A1;
14'd2565:data <=32'hFFB800B2;14'd2566:data <=32'hFFD300BD;14'd2567:data <=32'hFFF300C2;
14'd2568:data <=32'h001300BE;14'd2569:data <=32'h002F00B3;14'd2570:data <=32'h004600A4;
14'd2571:data <=32'h00590092;14'd2572:data <=32'h0069007E;14'd2573:data <=32'h00750069;
14'd2574:data <=32'h007C0052;14'd2575:data <=32'h007F003B;14'd2576:data <=32'h007C0023;
14'd2577:data <=32'h0072000E;14'd2578:data <=32'h0062FFFF;14'd2579:data <=32'h0051FFF6;
14'd2580:data <=32'h0040FFF7;14'd2581:data <=32'h0034FFFE;14'd2582:data <=32'h00310008;
14'd2583:data <=32'h00340012;14'd2584:data <=32'h003E0018;14'd2585:data <=32'h004B0015;
14'd2586:data <=32'h0056000C;14'd2587:data <=32'h005DFFFF;14'd2588:data <=32'h005EFFEF;
14'd2589:data <=32'h005AFFDE;14'd2590:data <=32'h0051FFD1;14'd2591:data <=32'h0046FFC8;
14'd2592:data <=32'h0038FFC3;14'd2593:data <=32'h002BFFC0;14'd2594:data <=32'h001EFFC3;
14'd2595:data <=32'h0012FFC7;14'd2596:data <=32'h0008FFD0;14'd2597:data <=32'h0000FFDC;
14'd2598:data <=32'hFFFFFFEA;14'd2599:data <=32'h0003FFFA;14'd2600:data <=32'h000F0007;
14'd2601:data <=32'h0023000F;14'd2602:data <=32'h003A000F;14'd2603:data <=32'h00520004;
14'd2604:data <=32'h0065FFF1;14'd2605:data <=32'h0071FFD4;14'd2606:data <=32'h0073FFB5;
14'd2607:data <=32'h006AFF96;14'd2608:data <=32'h0059FF7B;14'd2609:data <=32'h0042FF66;
14'd2610:data <=32'h0028FF58;14'd2611:data <=32'h000DFF50;14'd2612:data <=32'hFFF2FF4D;
14'd2613:data <=32'hFFD9FF4C;14'd2614:data <=32'hFFBFFF50;14'd2615:data <=32'hFFA5FF57;
14'd2616:data <=32'hFF8CFF62;14'd2617:data <=32'hFF74FF72;14'd2618:data <=32'hFF61FF86;
14'd2619:data <=32'hFF51FF9D;14'd2620:data <=32'hFF46FFB4;14'd2621:data <=32'hFF40FFCB;
14'd2622:data <=32'hFF39FFE1;14'd2623:data <=32'hFF34FFF5;14'd2624:data <=32'hFF9C0055;
14'd2625:data <=32'hFFA20051;14'd2626:data <=32'hFF950048;14'd2627:data <=32'hFF14002E;
14'd2628:data <=32'hFEE10046;14'd2629:data <=32'hFEF10080;14'd2630:data <=32'hFF1000B4;
14'd2631:data <=32'hFF3C00DF;14'd2632:data <=32'hFF7100FA;14'd2633:data <=32'hFFAA0107;
14'd2634:data <=32'hFFDF0105;14'd2635:data <=32'h001000F8;14'd2636:data <=32'h003A00E3;
14'd2637:data <=32'h005D00C5;14'd2638:data <=32'h007700A2;14'd2639:data <=32'h0087007C;
14'd2640:data <=32'h008D0053;14'd2641:data <=32'h0087002D;14'd2642:data <=32'h0076000B;
14'd2643:data <=32'h005CFFF4;14'd2644:data <=32'h003FFFE9;14'd2645:data <=32'h0023FFEB;
14'd2646:data <=32'h000DFFF7;14'd2647:data <=32'h00010009;14'd2648:data <=32'hFFFF001B;
14'd2649:data <=32'h0004002B;14'd2650:data <=32'h000F0036;14'd2651:data <=32'h001D003B;
14'd2652:data <=32'h0028003A;14'd2653:data <=32'h00330036;14'd2654:data <=32'h003B0030;
14'd2655:data <=32'h0041002A;14'd2656:data <=32'h00470024;14'd2657:data <=32'h004C001C;
14'd2658:data <=32'h004E0013;14'd2659:data <=32'h0050000A;14'd2660:data <=32'h004E0001;
14'd2661:data <=32'h004BFFFA;14'd2662:data <=32'h0046FFF5;14'd2663:data <=32'h0042FFF3;
14'd2664:data <=32'h003FFFF4;14'd2665:data <=32'h0040FFF4;14'd2666:data <=32'h0044FFF5;
14'd2667:data <=32'h004AFFF1;14'd2668:data <=32'h0050FFE9;14'd2669:data <=32'h0053FFDF;
14'd2670:data <=32'h0052FFD1;14'd2671:data <=32'h004CFFC6;14'd2672:data <=32'h0043FFBD;
14'd2673:data <=32'h003AFFBB;14'd2674:data <=32'h0033FFBC;14'd2675:data <=32'h0030FFBD;
14'd2676:data <=32'h0033FFBE;14'd2677:data <=32'h0038FFBB;14'd2678:data <=32'h0040FFB2;
14'd2679:data <=32'h0043FFA3;14'd2680:data <=32'h0043FF90;14'd2681:data <=32'h003DFF7A;
14'd2682:data <=32'h0031FF64;14'd2683:data <=32'h001EFF50;14'd2684:data <=32'h0006FF3E;
14'd2685:data <=32'hFFE8FF2F;14'd2686:data <=32'hFFC4FF24;14'd2687:data <=32'hFF9BFF1F;
14'd2688:data <=32'hFF7AFFBD;14'd2689:data <=32'hFF6DFFBE;14'd2690:data <=32'hFF6CFFB3;
14'd2691:data <=32'hFF5DFF45;14'd2692:data <=32'hFEFCFF4F;14'd2693:data <=32'hFED9FF89;
14'd2694:data <=32'hFEC9FFC8;14'd2695:data <=32'hFECA000A;14'd2696:data <=32'hFEDB0046;
14'd2697:data <=32'hFEF90078;14'd2698:data <=32'hFF1E009E;14'd2699:data <=32'hFF4700BB;
14'd2700:data <=32'hFF7500CE;14'd2701:data <=32'hFFA000D7;14'd2702:data <=32'hFFCD00D6;
14'd2703:data <=32'hFFF600CC;14'd2704:data <=32'h001900B8;14'd2705:data <=32'h0033009E;
14'd2706:data <=32'h0046007F;14'd2707:data <=32'h004C0060;14'd2708:data <=32'h00480046;
14'd2709:data <=32'h003E0032;14'd2710:data <=32'h00330026;14'd2711:data <=32'h00290021;
14'd2712:data <=32'h0022001F;14'd2713:data <=32'h001E001E;14'd2714:data <=32'h001C001C;
14'd2715:data <=32'h00190017;14'd2716:data <=32'h00130014;14'd2717:data <=32'h000C0011;
14'd2718:data <=32'h00030014;14'd2719:data <=32'hFFFB001A;14'd2720:data <=32'hFFF50024;
14'd2721:data <=32'hFFF40031;14'd2722:data <=32'hFFF7003F;14'd2723:data <=32'h0001004B;
14'd2724:data <=32'h000D0054;14'd2725:data <=32'h001C0059;14'd2726:data <=32'h002C005C;
14'd2727:data <=32'h003D005B;14'd2728:data <=32'h004E0057;14'd2729:data <=32'h005F004F;
14'd2730:data <=32'h00710042;14'd2731:data <=32'h00800032;14'd2732:data <=32'h008A001B;
14'd2733:data <=32'h008E0001;14'd2734:data <=32'h008BFFE6;14'd2735:data <=32'h007EFFCE;
14'd2736:data <=32'h006AFFBC;14'd2737:data <=32'h0054FFB5;14'd2738:data <=32'h003EFFB6;
14'd2739:data <=32'h002DFFC0;14'd2740:data <=32'h0025FFCE;14'd2741:data <=32'h0026FFDD;
14'd2742:data <=32'h002FFFE8;14'd2743:data <=32'h003EFFEC;14'd2744:data <=32'h004FFFE8;
14'd2745:data <=32'h005FFFDD;14'd2746:data <=32'h006CFFCB;14'd2747:data <=32'h0074FFB4;
14'd2748:data <=32'h0078FF99;14'd2749:data <=32'h0074FF7A;14'd2750:data <=32'h0067FF59;
14'd2751:data <=32'h0051FF37;14'd2752:data <=32'h0036FF61;14'd2753:data <=32'h0021FF39;
14'd2754:data <=32'h000DFF29;14'd2755:data <=32'h0013FF3F;14'd2756:data <=32'hFFB7FF20;
14'd2757:data <=32'hFF8FFF33;14'd2758:data <=32'hFF6FFF4E;14'd2759:data <=32'hFF58FF6F;
14'd2760:data <=32'hFF4BFF90;14'd2761:data <=32'hFF47FFAF;14'd2762:data <=32'hFF46FFCA;
14'd2763:data <=32'hFF48FFE2;14'd2764:data <=32'hFF4BFFF8;14'd2765:data <=32'hFF4F000E;
14'd2766:data <=32'hFF560023;14'd2767:data <=32'hFF610039;14'd2768:data <=32'hFF6F004B;
14'd2769:data <=32'hFF7F0059;14'd2770:data <=32'hFF910063;14'd2771:data <=32'hFFA0006A;
14'd2772:data <=32'hFFB00070;14'd2773:data <=32'hFFBF0076;14'd2774:data <=32'hFFCE007B;
14'd2775:data <=32'hFFE1007F;14'd2776:data <=32'hFFF6007F;14'd2777:data <=32'h000F007A;
14'd2778:data <=32'h0025006C;14'd2779:data <=32'h00370058;14'd2780:data <=32'h0041003E;
14'd2781:data <=32'h00410022;14'd2782:data <=32'h00360009;14'd2783:data <=32'h0024FFF6;
14'd2784:data <=32'h000CFFED;14'd2785:data <=32'hFFF5FFED;14'd2786:data <=32'hFFDFFFF6;
14'd2787:data <=32'hFFCE0005;14'd2788:data <=32'hFFC30017;14'd2789:data <=32'hFFBE002D;
14'd2790:data <=32'hFFBF0045;14'd2791:data <=32'hFFC6005C;14'd2792:data <=32'hFFD40071;
14'd2793:data <=32'hFFE80084;14'd2794:data <=32'h00030090;14'd2795:data <=32'h00200096;
14'd2796:data <=32'h00400093;14'd2797:data <=32'h005F0085;14'd2798:data <=32'h00760071;
14'd2799:data <=32'h00850056;14'd2800:data <=32'h008C003C;14'd2801:data <=32'h008A0024;
14'd2802:data <=32'h00840012;14'd2803:data <=32'h007A0007;14'd2804:data <=32'h00740001;
14'd2805:data <=32'h0072FFFF;14'd2806:data <=32'h0074FFFD;14'd2807:data <=32'h0079FFF6;
14'd2808:data <=32'h007FFFED;14'd2809:data <=32'h0083FFDF;14'd2810:data <=32'h0086FFCF;
14'd2811:data <=32'h0085FFBD;14'd2812:data <=32'h0081FFAC;14'd2813:data <=32'h007CFF9A;
14'd2814:data <=32'h0074FF88;14'd2815:data <=32'h0069FF74;14'd2816:data <=32'h00B1FFF4;
14'd2817:data <=32'h00CCFFBA;14'd2818:data <=32'h00C1FF81;14'd2819:data <=32'h0036FF6E;
14'd2820:data <=32'hFFE9FF51;14'd2821:data <=32'hFFD1FF65;14'd2822:data <=32'hFFC1FF7C;
14'd2823:data <=32'hFFBAFF94;14'd2824:data <=32'hFFBEFFA9;14'd2825:data <=32'hFFC6FFB6;
14'd2826:data <=32'hFFD0FFBA;14'd2827:data <=32'hFFD8FFB5;14'd2828:data <=32'hFFD8FFAE;
14'd2829:data <=32'hFFD2FFA4;14'd2830:data <=32'hFFC6FF9F;14'd2831:data <=32'hFFB4FF9D;
14'd2832:data <=32'hFFA4FFA0;14'd2833:data <=32'hFF92FFA7;14'd2834:data <=32'hFF81FFB4;
14'd2835:data <=32'hFF70FFC4;14'd2836:data <=32'hFF62FFD9;14'd2837:data <=32'hFF58FFF3;
14'd2838:data <=32'hFF540012;14'd2839:data <=32'hFF590035;14'd2840:data <=32'hFF680055;
14'd2841:data <=32'hFF820071;14'd2842:data <=32'hFFA40083;14'd2843:data <=32'hFFC90089;
14'd2844:data <=32'hFFEC0083;14'd2845:data <=32'h000A0072;14'd2846:data <=32'h001E005A;
14'd2847:data <=32'h0028003F;14'd2848:data <=32'h00280026;14'd2849:data <=32'h00210011;
14'd2850:data <=32'h00140001;14'd2851:data <=32'h0006FFF6;14'd2852:data <=32'hFFF6FFF1;
14'd2853:data <=32'hFFE4FFEF;14'd2854:data <=32'hFFD3FFF3;14'd2855:data <=32'hFFC4FFFC;
14'd2856:data <=32'hFFB60009;14'd2857:data <=32'hFFAB001C;14'd2858:data <=32'hFFA60032;
14'd2859:data <=32'hFFA70049;14'd2860:data <=32'hFFB0005F;14'd2861:data <=32'hFFBC0072;
14'd2862:data <=32'hFFCD0081;14'd2863:data <=32'hFFDF008C;14'd2864:data <=32'hFFF10093;
14'd2865:data <=32'h00020099;14'd2866:data <=32'h0014009F;14'd2867:data <=32'h002700A5;
14'd2868:data <=32'h004000AC;14'd2869:data <=32'h005D00AD;14'd2870:data <=32'h007F00A8;
14'd2871:data <=32'h00A3009A;14'd2872:data <=32'h00C50081;14'd2873:data <=32'h00E1005E;
14'd2874:data <=32'h00F30034;14'd2875:data <=32'h00FA0007;14'd2876:data <=32'h00F7FFDB;
14'd2877:data <=32'h00EBFFB0;14'd2878:data <=32'h00D7FF8B;14'd2879:data <=32'h00BBFF6A;
14'd2880:data <=32'h0071004B;14'd2881:data <=32'h00A50035;14'd2882:data <=32'h00CAFFFD;
14'd2883:data <=32'h0094FF54;14'd2884:data <=32'h0037FF2D;14'd2885:data <=32'h000BFF3B;
14'd2886:data <=32'hFFE9FF55;14'd2887:data <=32'hFFD2FF74;14'd2888:data <=32'hFFCAFF96;
14'd2889:data <=32'hFFD1FFB3;14'd2890:data <=32'hFFDEFFC6;14'd2891:data <=32'hFFEEFFCD;
14'd2892:data <=32'hFFFDFFCC;14'd2893:data <=32'h0007FFC4;14'd2894:data <=32'h000AFFB9;
14'd2895:data <=32'h0008FFAC;14'd2896:data <=32'h0001FFA2;14'd2897:data <=32'hFFF6FF98;
14'd2898:data <=32'hFFE8FF90;14'd2899:data <=32'hFFD7FF8D;14'd2900:data <=32'hFFC3FF8C;
14'd2901:data <=32'hFFADFF91;14'd2902:data <=32'hFF96FF9E;14'd2903:data <=32'hFF83FFB1;
14'd2904:data <=32'hFF77FFCC;14'd2905:data <=32'hFF73FFE8;14'd2906:data <=32'hFF790004;
14'd2907:data <=32'hFF87001A;14'd2908:data <=32'hFF98002A;14'd2909:data <=32'hFFAC0032;
14'd2910:data <=32'hFFBC0033;14'd2911:data <=32'hFFC90031;14'd2912:data <=32'hFFD3002E;
14'd2913:data <=32'hFFD8002B;14'd2914:data <=32'hFFDE0029;14'd2915:data <=32'hFFE50027;
14'd2916:data <=32'hFFEB0022;14'd2917:data <=32'hFFF1001D;14'd2918:data <=32'hFFF40015;
14'd2919:data <=32'hFFF5000A;14'd2920:data <=32'hFFF2FFFF;14'd2921:data <=32'hFFE9FFF5;
14'd2922:data <=32'hFFDEFFF0;14'd2923:data <=32'hFFCFFFED;14'd2924:data <=32'hFFC1FFEF;
14'd2925:data <=32'hFFB1FFF4;14'd2926:data <=32'hFFA1FFFD;14'd2927:data <=32'hFF92000A;
14'd2928:data <=32'hFF83001C;14'd2929:data <=32'hFF760035;14'd2930:data <=32'hFF6C0055;
14'd2931:data <=32'hFF6C007B;14'd2932:data <=32'hFF7600A6;14'd2933:data <=32'hFF8E00D0;
14'd2934:data <=32'hFFB400F8;14'd2935:data <=32'hFFE90113;14'd2936:data <=32'h00230120;
14'd2937:data <=32'h0062011C;14'd2938:data <=32'h009D0106;14'd2939:data <=32'h00D000E2;
14'd2940:data <=32'h00F800B6;14'd2941:data <=32'h01140080;14'd2942:data <=32'h0123004A;
14'd2943:data <=32'h01270012;14'd2944:data <=32'h00820050;14'd2945:data <=32'h00A70045;
14'd2946:data <=32'h00D50033;14'd2947:data <=32'h011DFFF4;14'd2948:data <=32'h00D6FFA6;
14'd2949:data <=32'h00B4FF8D;14'd2950:data <=32'h0092FF80;14'd2951:data <=32'h0073FF7C;
14'd2952:data <=32'h005AFF81;14'd2953:data <=32'h004BFF88;14'd2954:data <=32'h0041FF8E;
14'd2955:data <=32'h003AFF8F;14'd2956:data <=32'h0032FF8D;14'd2957:data <=32'h0029FF88;
14'd2958:data <=32'h001CFF86;14'd2959:data <=32'h000DFF85;14'd2960:data <=32'hFFFEFF89;
14'd2961:data <=32'hFFF2FF8F;14'd2962:data <=32'hFFE6FF97;14'd2963:data <=32'hFFDFFF9F;
14'd2964:data <=32'hFFD8FFA7;14'd2965:data <=32'hFFD3FFAE;14'd2966:data <=32'hFFCDFFB6;
14'd2967:data <=32'hFFC8FFBF;14'd2968:data <=32'hFFC6FFCB;14'd2969:data <=32'hFFC6FFD5;
14'd2970:data <=32'hFFCCFFDF;14'd2971:data <=32'hFFD4FFE4;14'd2972:data <=32'hFFDDFFE6;
14'd2973:data <=32'hFFE2FFE0;14'd2974:data <=32'hFFE3FFD9;14'd2975:data <=32'hFFDEFFD0;
14'd2976:data <=32'hFFD5FFCB;14'd2977:data <=32'hFFC8FFCC;14'd2978:data <=32'hFFBBFFD2;
14'd2979:data <=32'hFFB1FFDE;14'd2980:data <=32'hFFAEFFED;14'd2981:data <=32'hFFB0FFFC;
14'd2982:data <=32'hFFB70008;14'd2983:data <=32'hFFC20010;14'd2984:data <=32'hFFCD0011;
14'd2985:data <=32'hFFD7000F;14'd2986:data <=32'hFFDF0009;14'd2987:data <=32'hFFE30001;
14'd2988:data <=32'hFFE3FFF6;14'd2989:data <=32'hFFDFFFEB;14'd2990:data <=32'hFFD6FFE1;
14'd2991:data <=32'hFFC9FFD7;14'd2992:data <=32'hFFB6FFD2;14'd2993:data <=32'hFF9CFFD3;
14'd2994:data <=32'hFF80FFDC;14'd2995:data <=32'hFF64FFF1;14'd2996:data <=32'hFF4D0011;
14'd2997:data <=32'hFF3F003A;14'd2998:data <=32'hFF400069;14'd2999:data <=32'hFF4E009A;
14'd3000:data <=32'hFF6B00C3;14'd3001:data <=32'hFF9200E4;14'd3002:data <=32'hFFBF00F8;
14'd3003:data <=32'hFFEE0100;14'd3004:data <=32'h001B00FF;14'd3005:data <=32'h004500F6;
14'd3006:data <=32'h006B00E5;14'd3007:data <=32'h008D00CF;14'd3008:data <=32'h007B00DB;
14'd3009:data <=32'h00AF00D0;14'd3010:data <=32'h00CF00C2;14'd3011:data <=32'h00A000CC;
14'd3012:data <=32'h0089008D;14'd3013:data <=32'h0097007C;14'd3014:data <=32'h00A2006A;
14'd3015:data <=32'h00AE0059;14'd3016:data <=32'h00BA0047;14'd3017:data <=32'h00C80033;
14'd3018:data <=32'h00D50018;14'd3019:data <=32'h00DFFFF6;14'd3020:data <=32'h00E0FFCF;
14'd3021:data <=32'h00D6FFA5;14'd3022:data <=32'h00C0FF7E;14'd3023:data <=32'h009FFF5E;
14'd3024:data <=32'h0077FF49;14'd3025:data <=32'h004DFF40;14'd3026:data <=32'h0024FF43;
14'd3027:data <=32'h0000FF4E;14'd3028:data <=32'hFFE2FF60;14'd3029:data <=32'hFFCAFF76;
14'd3030:data <=32'hFFBAFF90;14'd3031:data <=32'hFFB0FFAC;14'd3032:data <=32'hFFAEFFC9;
14'd3033:data <=32'hFFB4FFE5;14'd3034:data <=32'hFFC3FFFD;14'd3035:data <=32'hFFD8000D;
14'd3036:data <=32'hFFF10014;14'd3037:data <=32'h000C000F;14'd3038:data <=32'h001F0001;
14'd3039:data <=32'h002BFFED;14'd3040:data <=32'h002EFFD6;14'd3041:data <=32'h0027FFC1;
14'd3042:data <=32'h001AFFB2;14'd3043:data <=32'h0008FFA9;14'd3044:data <=32'hFFF8FFA6;
14'd3045:data <=32'hFFEAFFA8;14'd3046:data <=32'hFFDEFFAD;14'd3047:data <=32'hFFD7FFB3;
14'd3048:data <=32'hFFD0FFB8;14'd3049:data <=32'hFFCAFFBC;14'd3050:data <=32'hFFC5FFC0;
14'd3051:data <=32'hFFBFFFC3;14'd3052:data <=32'hFFBBFFC8;14'd3053:data <=32'hFFB6FFCC;
14'd3054:data <=32'hFFB2FFD0;14'd3055:data <=32'hFFAEFFD2;14'd3056:data <=32'hFFA8FFD4;
14'd3057:data <=32'hFF9FFFD5;14'd3058:data <=32'hFF93FFDA;14'd3059:data <=32'hFF85FFE2;
14'd3060:data <=32'hFF75FFF1;14'd3061:data <=32'hFF6B0005;14'd3062:data <=32'hFF66001F;
14'd3063:data <=32'hFF68003A;14'd3064:data <=32'hFF730054;14'd3065:data <=32'hFF830067;
14'd3066:data <=32'hFF960074;14'd3067:data <=32'hFFA8007A;14'd3068:data <=32'hFFB6007D;
14'd3069:data <=32'hFFC2007F;14'd3070:data <=32'hFFCA0082;14'd3071:data <=32'hFFD00088;
14'd3072:data <=32'hFFAC0109;14'd3073:data <=32'hFFE10129;14'd3074:data <=32'h00110123;
14'd3075:data <=32'hFFDD00A7;14'd3076:data <=32'hFFBC008D;14'd3077:data <=32'hFFC800A3;
14'd3078:data <=32'hFFDB00B9;14'd3079:data <=32'hFFF500CC;14'd3080:data <=32'h001700DD;
14'd3081:data <=32'h004100E6;14'd3082:data <=32'h007200E4;14'd3083:data <=32'h00A500D1;
14'd3084:data <=32'h00D300B0;14'd3085:data <=32'h00F60081;14'd3086:data <=32'h010B0049;
14'd3087:data <=32'h010E000F;14'd3088:data <=32'h0101FFD8;14'd3089:data <=32'h00E9FFA9;
14'd3090:data <=32'h00C8FF85;14'd3091:data <=32'h00A1FF6C;14'd3092:data <=32'h0079FF5B;
14'd3093:data <=32'h0050FF56;14'd3094:data <=32'h0029FF58;14'd3095:data <=32'h0005FF65;
14'd3096:data <=32'hFFE6FF78;14'd3097:data <=32'hFFCFFF93;14'd3098:data <=32'hFFC3FFB2;
14'd3099:data <=32'hFFC1FFD1;14'd3100:data <=32'hFFC9FFEE;14'd3101:data <=32'hFFD90002;
14'd3102:data <=32'hFFEE0010;14'd3103:data <=32'h00020013;14'd3104:data <=32'h00140011;
14'd3105:data <=32'h0022000A;14'd3106:data <=32'h002C0001;14'd3107:data <=32'h0033FFF7;
14'd3108:data <=32'h0038FFEF;14'd3109:data <=32'h003FFFE4;14'd3110:data <=32'h0045FFD9;
14'd3111:data <=32'h0049FFCA;14'd3112:data <=32'h004AFFB7;14'd3113:data <=32'h0047FFA2;
14'd3114:data <=32'h003DFF8C;14'd3115:data <=32'h002CFF78;14'd3116:data <=32'h0016FF68;
14'd3117:data <=32'hFFFBFF5E;14'd3118:data <=32'hFFDEFF5A;14'd3119:data <=32'hFFC1FF5C;
14'd3120:data <=32'hFFA5FF63;14'd3121:data <=32'hFF8AFF70;14'd3122:data <=32'hFF71FF83;
14'd3123:data <=32'hFF5BFF9A;14'd3124:data <=32'hFF48FFB7;14'd3125:data <=32'hFF3DFFD9;
14'd3126:data <=32'hFF3DFFFF;14'd3127:data <=32'hFF460023;14'd3128:data <=32'hFF590042;
14'd3129:data <=32'hFF750058;14'd3130:data <=32'hFF930062;14'd3131:data <=32'hFFB00061;
14'd3132:data <=32'hFFC50057;14'd3133:data <=32'hFFD10047;14'd3134:data <=32'hFFD30039;
14'd3135:data <=32'hFFCD002D;14'd3136:data <=32'hFF490054;14'd3137:data <=32'hFF4A007F;
14'd3138:data <=32'hFF6E009E;14'd3139:data <=32'hFFC70059;14'd3140:data <=32'hFF970035;
14'd3141:data <=32'hFF8F0046;14'd3142:data <=32'hFF8B005D;14'd3143:data <=32'hFF8D0077;
14'd3144:data <=32'hFF970095;14'd3145:data <=32'hFFAC00B3;14'd3146:data <=32'hFFCB00CC;
14'd3147:data <=32'hFFF300DD;14'd3148:data <=32'h002200E0;14'd3149:data <=32'h004E00D5;
14'd3150:data <=32'h007500BF;14'd3151:data <=32'h0092009F;14'd3152:data <=32'h00A5007C;
14'd3153:data <=32'h00AE005A;14'd3154:data <=32'h00AF003A;14'd3155:data <=32'h00AB001D;
14'd3156:data <=32'h00A40005;14'd3157:data <=32'h009AFFEE;14'd3158:data <=32'h008DFFD8;
14'd3159:data <=32'h007DFFC7;14'd3160:data <=32'h006AFFBA;14'd3161:data <=32'h0053FFB2;
14'd3162:data <=32'h003EFFB0;14'd3163:data <=32'h002BFFB4;14'd3164:data <=32'h001DFFBA;
14'd3165:data <=32'h0011FFC4;14'd3166:data <=32'h000BFFCC;14'd3167:data <=32'h0004FFD5;
14'd3168:data <=32'h0000FFDD;14'd3169:data <=32'hFFFBFFE6;14'd3170:data <=32'hFFF7FFF2;
14'd3171:data <=32'hFFF80000;14'd3172:data <=32'hFFFC0011;14'd3173:data <=32'h00090021;
14'd3174:data <=32'h001D002E;14'd3175:data <=32'h00380032;14'd3176:data <=32'h0056002D;
14'd3177:data <=32'h0072001D;14'd3178:data <=32'h00880002;14'd3179:data <=32'h0097FFE0;
14'd3180:data <=32'h009CFFBA;14'd3181:data <=32'h0095FF93;14'd3182:data <=32'h0084FF6E;
14'd3183:data <=32'h006BFF4F;14'd3184:data <=32'h004BFF35;14'd3185:data <=32'h0025FF23;
14'd3186:data <=32'hFFFAFF19;14'd3187:data <=32'hFFCDFF1A;14'd3188:data <=32'hFFA1FF25;
14'd3189:data <=32'hFF77FF3C;14'd3190:data <=32'hFF56FF5E;14'd3191:data <=32'hFF40FF86;
14'd3192:data <=32'hFF37FFB1;14'd3193:data <=32'hFF3BFFDB;14'd3194:data <=32'hFF4AFFFC;
14'd3195:data <=32'hFF5F0013;14'd3196:data <=32'hFF740020;14'd3197:data <=32'hFF850024;
14'd3198:data <=32'hFF920023;14'd3199:data <=32'hFF980020;14'd3200:data <=32'hFFA4FFFB;
14'd3201:data <=32'hFF93FFFD;14'd3202:data <=32'hFF870016;14'd3203:data <=32'hFF800058;
14'd3204:data <=32'hFF62003A;14'd3205:data <=32'hFF69004D;14'd3206:data <=32'hFF73005F;
14'd3207:data <=32'hFF7F006F;14'd3208:data <=32'hFF8D0080;14'd3209:data <=32'hFFA00090;
14'd3210:data <=32'hFFB8009F;14'd3211:data <=32'hFFD300A6;14'd3212:data <=32'hFFF100A7;
14'd3213:data <=32'h000E009E;14'd3214:data <=32'h0024008C;14'd3215:data <=32'h00330078;
14'd3216:data <=32'h00390063;14'd3217:data <=32'h00360052;14'd3218:data <=32'h00310047;
14'd3219:data <=32'h002B0043;14'd3220:data <=32'h00290044;14'd3221:data <=32'h002B0045;
14'd3222:data <=32'h00300047;14'd3223:data <=32'h00380046;14'd3224:data <=32'h00410042;
14'd3225:data <=32'h004A003C;14'd3226:data <=32'h00500033;14'd3227:data <=32'h00560029;
14'd3228:data <=32'h005B001F;14'd3229:data <=32'h005E0012;14'd3230:data <=32'h005E0004;
14'd3231:data <=32'h005BFFF4;14'd3232:data <=32'h0051FFE4;14'd3233:data <=32'h0043FFD8;
14'd3234:data <=32'h002FFFD1;14'd3235:data <=32'h0019FFD3;14'd3236:data <=32'h0006FFDE;
14'd3237:data <=32'hFFF8FFF0;14'd3238:data <=32'hFFF50008;14'd3239:data <=32'hFFFB0020;
14'd3240:data <=32'h000A0033;14'd3241:data <=32'h00230041;14'd3242:data <=32'h003E0044;
14'd3243:data <=32'h0059003E;14'd3244:data <=32'h00720030;14'd3245:data <=32'h0086001C;
14'd3246:data <=32'h00950002;14'd3247:data <=32'h009DFFE7;14'd3248:data <=32'h00A0FFCA;
14'd3249:data <=32'h009DFFAA;14'd3250:data <=32'h0094FF8B;14'd3251:data <=32'h0082FF6E;
14'd3252:data <=32'h0069FF56;14'd3253:data <=32'h004DFF43;14'd3254:data <=32'h002BFF39;
14'd3255:data <=32'h000AFF37;14'd3256:data <=32'hFFEDFF3C;14'd3257:data <=32'hFFD5FF44;
14'd3258:data <=32'hFFC2FF4F;14'd3259:data <=32'hFFB2FF58;14'd3260:data <=32'hFFA3FF5E;
14'd3261:data <=32'hFF91FF64;14'd3262:data <=32'hFF7CFF6B;14'd3263:data <=32'hFF63FF77;
14'd3264:data <=32'hFFA6FFFF;14'd3265:data <=32'hFFA8FFF6;14'd3266:data <=32'hFF9DFFE8;
14'd3267:data <=32'hFF29FFB0;14'd3268:data <=32'hFEF4FFAD;14'd3269:data <=32'hFEECFFE1;
14'd3270:data <=32'hFEF00012;14'd3271:data <=32'hFEFF0043;14'd3272:data <=32'hFF16006D;
14'd3273:data <=32'hFF350092;14'd3274:data <=32'hFF5B00AF;14'd3275:data <=32'hFF8900C2;
14'd3276:data <=32'hFFB900C8;14'd3277:data <=32'hFFE700BF;14'd3278:data <=32'h000F00AB;
14'd3279:data <=32'h002B008B;14'd3280:data <=32'h00390068;14'd3281:data <=32'h00390047;
14'd3282:data <=32'h002E002C;14'd3283:data <=32'h001E001C;14'd3284:data <=32'h000C0015;
14'd3285:data <=32'hFFFC0017;14'd3286:data <=32'hFFF0001E;14'd3287:data <=32'hFFEA0028;
14'd3288:data <=32'hFFE80033;14'd3289:data <=32'hFFEA003E;14'd3290:data <=32'hFFEF0048;
14'd3291:data <=32'hFFF70051;14'd3292:data <=32'h00030058;14'd3293:data <=32'h0012005C;
14'd3294:data <=32'h0022005B;14'd3295:data <=32'h00320055;14'd3296:data <=32'h003F0048;
14'd3297:data <=32'h00460039;14'd3298:data <=32'h0048002A;14'd3299:data <=32'h0043001B;
14'd3300:data <=32'h003A0012;14'd3301:data <=32'h002F000F;14'd3302:data <=32'h00280012;
14'd3303:data <=32'h00230018;14'd3304:data <=32'h00250020;14'd3305:data <=32'h002B0026;
14'd3306:data <=32'h00320028;14'd3307:data <=32'h003A0027;14'd3308:data <=32'h00420023;
14'd3309:data <=32'h0047001E;14'd3310:data <=32'h004A0019;14'd3311:data <=32'h004D0016;
14'd3312:data <=32'h00510014;14'd3313:data <=32'h00580012;14'd3314:data <=32'h0060000E;
14'd3315:data <=32'h006A0008;14'd3316:data <=32'h0074FFFF;14'd3317:data <=32'h007CFFF2;
14'd3318:data <=32'h0084FFE5;14'd3319:data <=32'h0089FFD4;14'd3320:data <=32'h008EFFC3;
14'd3321:data <=32'h0092FFAD;14'd3322:data <=32'h0096FF93;14'd3323:data <=32'h0095FF75;
14'd3324:data <=32'h008BFF50;14'd3325:data <=32'h0077FF2A;14'd3326:data <=32'h0055FF05;
14'd3327:data <=32'h0026FEE9;14'd3328:data <=32'hFFC4FF8B;14'd3329:data <=32'hFFBBFF84;
14'd3330:data <=32'hFFC0FF75;14'd3331:data <=32'hFFD1FEFE;14'd3332:data <=32'hFF77FEE0;
14'd3333:data <=32'hFF43FF03;14'd3334:data <=32'hFF1AFF2F;14'd3335:data <=32'hFEFDFF63;
14'd3336:data <=32'hFEEBFF9A;14'd3337:data <=32'hFEE6FFD2;14'd3338:data <=32'hFEEE000A;
14'd3339:data <=32'hFF03003D;14'd3340:data <=32'hFF240068;14'd3341:data <=32'hFF4E0085;
14'd3342:data <=32'hFF7C0094;14'd3343:data <=32'hFFA70096;14'd3344:data <=32'hFFCB008A;
14'd3345:data <=32'hFFE50079;14'd3346:data <=32'hFFF50065;14'd3347:data <=32'hFFFB0053;
14'd3348:data <=32'hFFFD0045;14'd3349:data <=32'hFFFD003B;14'd3350:data <=32'hFFFC0033;
14'd3351:data <=32'hFFFD002E;14'd3352:data <=32'hFFFC0028;14'd3353:data <=32'hFFFB0022;
14'd3354:data <=32'hFFF5001E;14'd3355:data <=32'hFFF0001C;14'd3356:data <=32'hFFEA001C;
14'd3357:data <=32'hFFE40021;14'd3358:data <=32'hFFE10027;14'd3359:data <=32'hFFE1002E;
14'd3360:data <=32'hFFE30034;14'd3361:data <=32'hFFE50039;14'd3362:data <=32'hFFE7003D;
14'd3363:data <=32'hFFE80041;14'd3364:data <=32'hFFE90049;14'd3365:data <=32'hFFED0052;
14'd3366:data <=32'hFFF5005D;14'd3367:data <=32'h00010067;14'd3368:data <=32'h0012006E;
14'd3369:data <=32'h00270070;14'd3370:data <=32'h003D006A;14'd3371:data <=32'h0050005D;
14'd3372:data <=32'h005D004A;14'd3373:data <=32'h00630036;14'd3374:data <=32'h00600022;
14'd3375:data <=32'h00580013;14'd3376:data <=32'h004D000A;14'd3377:data <=32'h00400007;
14'd3378:data <=32'h0037000A;14'd3379:data <=32'h00320012;14'd3380:data <=32'h0031001B;
14'd3381:data <=32'h00350025;14'd3382:data <=32'h003D002E;14'd3383:data <=32'h004B0036;
14'd3384:data <=32'h005E003C;14'd3385:data <=32'h0077003C;14'd3386:data <=32'h00950034;
14'd3387:data <=32'h00B40020;14'd3388:data <=32'h00D00000;14'd3389:data <=32'h00E2FFD3;
14'd3390:data <=32'h00E9FF9E;14'd3391:data <=32'h00DEFF67;14'd3392:data <=32'h008CFF8A;
14'd3393:data <=32'h0089FF5F;14'd3394:data <=32'h0083FF4B;14'd3395:data <=32'h0092FF58;
14'd3396:data <=32'h004DFF13;14'd3397:data <=32'h0023FF0E;14'd3398:data <=32'hFFFCFF10;
14'd3399:data <=32'hFFD8FF19;14'd3400:data <=32'hFFB6FF27;14'd3401:data <=32'hFF97FF39;
14'd3402:data <=32'hFF7CFF52;14'd3403:data <=32'hFF69FF6F;14'd3404:data <=32'hFF5EFF8F;
14'd3405:data <=32'hFF58FFAD;14'd3406:data <=32'hFF5DFFC8;14'd3407:data <=32'hFF62FFDD;
14'd3408:data <=32'hFF69FFED;14'd3409:data <=32'hFF6DFFFC;14'd3410:data <=32'hFF720008;
14'd3411:data <=32'hFF740018;14'd3412:data <=32'hFF790029;14'd3413:data <=32'hFF83003D;
14'd3414:data <=32'hFF920050;14'd3415:data <=32'hFFA8005D;14'd3416:data <=32'hFFC00065;
14'd3417:data <=32'hFFDA0063;14'd3418:data <=32'hFFF1005A;14'd3419:data <=32'h0003004B;
14'd3420:data <=32'h000D0039;14'd3421:data <=32'h00110026;14'd3422:data <=32'h00100015;
14'd3423:data <=32'h000A0005;14'd3424:data <=32'h0000FFF9;14'd3425:data <=32'hFFF2FFF0;
14'd3426:data <=32'hFFE0FFEA;14'd3427:data <=32'hFFCCFFEB;14'd3428:data <=32'hFFB7FFF4;
14'd3429:data <=32'hFFA50003;14'd3430:data <=32'hFF98001C;14'd3431:data <=32'hFF930039;
14'd3432:data <=32'hFF990056;14'd3433:data <=32'hFFA90071;14'd3434:data <=32'hFFC20087;
14'd3435:data <=32'hFFDE0092;14'd3436:data <=32'hFFFB0094;14'd3437:data <=32'h0015008C;
14'd3438:data <=32'h00280080;14'd3439:data <=32'h00350072;14'd3440:data <=32'h003C0065;
14'd3441:data <=32'h003F005A;14'd3442:data <=32'h00410051;14'd3443:data <=32'h0043004C;
14'd3444:data <=32'h00440049;14'd3445:data <=32'h00470047;14'd3446:data <=32'h004B0045;
14'd3447:data <=32'h004F0046;14'd3448:data <=32'h00560047;14'd3449:data <=32'h00610048;
14'd3450:data <=32'h00700048;14'd3451:data <=32'h00850043;14'd3452:data <=32'h009A0037;
14'd3453:data <=32'h00B00022;14'd3454:data <=32'h00BF0004;14'd3455:data <=32'h00C7FFE0;
14'd3456:data <=32'h00C50057;14'd3457:data <=32'h00F4002C;14'd3458:data <=32'h00FFFFFA;
14'd3459:data <=32'h008EFFC4;14'd3460:data <=32'h005DFF8A;14'd3461:data <=32'h004AFF8C;
14'd3462:data <=32'h003DFF91;14'd3463:data <=32'h0036FF96;14'd3464:data <=32'h0032FF97;
14'd3465:data <=32'h002FFF94;14'd3466:data <=32'h002AFF91;14'd3467:data <=32'h0024FF8C;
14'd3468:data <=32'h001DFF85;14'd3469:data <=32'h0016FF7F;14'd3470:data <=32'h000CFF78;
14'd3471:data <=32'hFFFFFF6F;14'd3472:data <=32'hFFEEFF65;14'd3473:data <=32'hFFD6FF5D;
14'd3474:data <=32'hFFB8FF5D;14'd3475:data <=32'hFF96FF65;14'd3476:data <=32'hFF77FF79;
14'd3477:data <=32'hFF5CFF97;14'd3478:data <=32'hFF4CFFBD;14'd3479:data <=32'hFF49FFE6;
14'd3480:data <=32'hFF52000E;14'd3481:data <=32'hFF66002F;14'd3482:data <=32'hFF810046;
14'd3483:data <=32'hFF9E0054;14'd3484:data <=32'hFFBB0059;14'd3485:data <=32'hFFD70056;
14'd3486:data <=32'hFFEF004D;14'd3487:data <=32'h0002003E;14'd3488:data <=32'h0011002C;
14'd3489:data <=32'h00180016;14'd3490:data <=32'h0018FFFF;14'd3491:data <=32'h0010FFE9;
14'd3492:data <=32'h0000FFD5;14'd3493:data <=32'hFFEBFFCA;14'd3494:data <=32'hFFD1FFC6;
14'd3495:data <=32'hFFB7FFCC;14'd3496:data <=32'hFFA1FFDA;14'd3497:data <=32'hFF93FFEE;
14'd3498:data <=32'hFF8A0005;14'd3499:data <=32'hFF870019;14'd3500:data <=32'hFF8B002C;
14'd3501:data <=32'hFF8F003D;14'd3502:data <=32'hFF93004B;14'd3503:data <=32'hFF97005A;
14'd3504:data <=32'hFF9B006A;14'd3505:data <=32'hFFA2007D;14'd3506:data <=32'hFFAE0092;
14'd3507:data <=32'hFFBF00A6;14'd3508:data <=32'hFFD700B7;14'd3509:data <=32'hFFF500C3;
14'd3510:data <=32'h001400C8;14'd3511:data <=32'h003500C8;14'd3512:data <=32'h005500C1;
14'd3513:data <=32'h007200B5;14'd3514:data <=32'h008F00A4;14'd3515:data <=32'h00AA008E;
14'd3516:data <=32'h00C20071;14'd3517:data <=32'h00D4004F;14'd3518:data <=32'h00DE0028;
14'd3519:data <=32'h00DDFFFD;14'd3520:data <=32'h004400A4;14'd3521:data <=32'h007E00A6;
14'd3522:data <=32'h00B50085;14'd3523:data <=32'h00B6FFD6;14'd3524:data <=32'h0079FF94;
14'd3525:data <=32'h0058FF97;14'd3526:data <=32'h003FFFA3;14'd3527:data <=32'h0030FFB5;
14'd3528:data <=32'h0029FFC4;14'd3529:data <=32'h002AFFD1;14'd3530:data <=32'h002EFFD9;
14'd3531:data <=32'h0037FFDE;14'd3532:data <=32'h0041FFDE;14'd3533:data <=32'h004BFFD9;
14'd3534:data <=32'h0056FFCF;14'd3535:data <=32'h005EFFBE;14'd3536:data <=32'h0061FFA6;
14'd3537:data <=32'h005AFF8C;14'd3538:data <=32'h004AFF72;14'd3539:data <=32'h002FFF5D;
14'd3540:data <=32'h000DFF51;14'd3541:data <=32'hFFE8FF51;14'd3542:data <=32'hFFC6FF5C;
14'd3543:data <=32'hFFAAFF71;14'd3544:data <=32'hFF96FF8B;14'd3545:data <=32'hFF8CFFA6;
14'd3546:data <=32'hFF8AFFC1;14'd3547:data <=32'hFF8DFFD8;14'd3548:data <=32'hFF93FFEC;
14'd3549:data <=32'hFF9CFFFC;14'd3550:data <=32'hFFA7000A;14'd3551:data <=32'hFFB20014;
14'd3552:data <=32'hFFC2001B;14'd3553:data <=32'hFFD1001E;14'd3554:data <=32'hFFE2001D;
14'd3555:data <=32'hFFEF0016;14'd3556:data <=32'hFFF9000B;14'd3557:data <=32'hFFFFFFFF;
14'd3558:data <=32'hFFFFFFF1;14'd3559:data <=32'hFFFBFFE6;14'd3560:data <=32'hFFF6FFDC;
14'd3561:data <=32'hFFEFFFD4;14'd3562:data <=32'hFFE6FFCD;14'd3563:data <=32'hFFDCFFC5;
14'd3564:data <=32'hFFD0FFBD;14'd3565:data <=32'hFFBFFFB7;14'd3566:data <=32'hFFA8FFB2;
14'd3567:data <=32'hFF8BFFB5;14'd3568:data <=32'hFF6CFFC1;14'd3569:data <=32'hFF4EFFD9;
14'd3570:data <=32'hFF34FFFB;14'd3571:data <=32'hFF230027;14'd3572:data <=32'hFF200059;
14'd3573:data <=32'hFF2B008B;14'd3574:data <=32'hFF4200BB;14'd3575:data <=32'hFF6400E3;
14'd3576:data <=32'hFF900103;14'd3577:data <=32'hFFC10118;14'd3578:data <=32'hFFF70124;
14'd3579:data <=32'h002E0123;14'd3580:data <=32'h00660116;14'd3581:data <=32'h009A00FB;
14'd3582:data <=32'h00C600D3;14'd3583:data <=32'h00E700A1;14'd3584:data <=32'h002B008F;
14'd3585:data <=32'h004D009B;14'd3586:data <=32'h007C00A2;14'd3587:data <=32'h00DF007A;
14'd3588:data <=32'h00BC0020;14'd3589:data <=32'h00AB0008;14'd3590:data <=32'h009AFFF9;
14'd3591:data <=32'h008BFFF1;14'd3592:data <=32'h0080FFEA;14'd3593:data <=32'h0078FFE4;
14'd3594:data <=32'h0071FFDF;14'd3595:data <=32'h006AFFD9;14'd3596:data <=32'h0064FFD4;
14'd3597:data <=32'h005FFFD1;14'd3598:data <=32'h005BFFCD;14'd3599:data <=32'h0059FFC8;
14'd3600:data <=32'h0058FFC1;14'd3601:data <=32'h0055FFB6;14'd3602:data <=32'h004FFFAA;
14'd3603:data <=32'h0043FF9E;14'd3604:data <=32'h0032FF96;14'd3605:data <=32'h001FFF93;
14'd3606:data <=32'h000CFF97;14'd3607:data <=32'hFFFFFFA1;14'd3608:data <=32'hFFF7FFAD;
14'd3609:data <=32'hFFF4FFB7;14'd3610:data <=32'hFFF6FFBF;14'd3611:data <=32'hFFF8FFC1;
14'd3612:data <=32'hFFFAFFC0;14'd3613:data <=32'hFFF7FFBC;14'd3614:data <=32'hFFF2FFB9;
14'd3615:data <=32'hFFEAFFB8;14'd3616:data <=32'hFFE1FFBB;14'd3617:data <=32'hFFD9FFC1;
14'd3618:data <=32'hFFD4FFC9;14'd3619:data <=32'hFFD1FFD2;14'd3620:data <=32'hFFD0FFD9;
14'd3621:data <=32'hFFD1FFE1;14'd3622:data <=32'hFFD4FFE8;14'd3623:data <=32'hFFD9FFEE;
14'd3624:data <=32'hFFDFFFF3;14'd3625:data <=32'hFFE9FFF6;14'd3626:data <=32'hFFF5FFF4;
14'd3627:data <=32'h0001FFEB;14'd3628:data <=32'h000AFFDD;14'd3629:data <=32'h000EFFC8;
14'd3630:data <=32'h0008FFAE;14'd3631:data <=32'hFFF8FF95;14'd3632:data <=32'hFFDCFF80;
14'd3633:data <=32'hFFB7FF76;14'd3634:data <=32'hFF8DFF77;14'd3635:data <=32'hFF64FF86;
14'd3636:data <=32'hFF3FFFA2;14'd3637:data <=32'hFF23FFC8;14'd3638:data <=32'hFF11FFF4;
14'd3639:data <=32'hFF0A0023;14'd3640:data <=32'hFF0E0052;14'd3641:data <=32'hFF1C007F;
14'd3642:data <=32'hFF3300A9;14'd3643:data <=32'hFF5200CF;14'd3644:data <=32'hFF7A00EE;
14'd3645:data <=32'hFFA80102;14'd3646:data <=32'hFFDB010A;14'd3647:data <=32'h000C0105;
14'd3648:data <=32'hFFFC00E7;14'd3649:data <=32'h002600F0;14'd3650:data <=32'h003F00F4;
14'd3651:data <=32'h001800FC;14'd3652:data <=32'h001700C0;14'd3653:data <=32'h002A00BF;
14'd3654:data <=32'h004000BE;14'd3655:data <=32'h005900BC;14'd3656:data <=32'h007600B3;
14'd3657:data <=32'h009400A2;14'd3658:data <=32'h00AF0088;14'd3659:data <=32'h00C30068;
14'd3660:data <=32'h00CF0044;14'd3661:data <=32'h00D2001F;14'd3662:data <=32'h00CDFFFB;
14'd3663:data <=32'h00C2FFDB;14'd3664:data <=32'h00B3FFBE;14'd3665:data <=32'h009DFFA6;
14'd3666:data <=32'h0083FF90;14'd3667:data <=32'h0064FF81;14'd3668:data <=32'h0042FF7B;
14'd3669:data <=32'h0020FF7F;14'd3670:data <=32'h0002FF8E;14'd3671:data <=32'hFFECFFA5;
14'd3672:data <=32'hFFE0FFC1;14'd3673:data <=32'hFFE1FFDD;14'd3674:data <=32'hFFEBFFF4;
14'd3675:data <=32'hFFFD0002;14'd3676:data <=32'h00100008;14'd3677:data <=32'h00230004;
14'd3678:data <=32'h0031FFFA;14'd3679:data <=32'h0038FFEC;14'd3680:data <=32'h003BFFDE;
14'd3681:data <=32'h0039FFD1;14'd3682:data <=32'h0034FFC5;14'd3683:data <=32'h002DFFBC;
14'd3684:data <=32'h0025FFB4;14'd3685:data <=32'h001AFFAE;14'd3686:data <=32'h000EFFAC;
14'd3687:data <=32'h0003FFAC;14'd3688:data <=32'hFFF9FFB0;14'd3689:data <=32'hFFF2FFB6;
14'd3690:data <=32'hFFEFFFBE;14'd3691:data <=32'hFFF1FFC4;14'd3692:data <=32'hFFF6FFC5;
14'd3693:data <=32'hFFFBFFC2;14'd3694:data <=32'h0000FFB9;14'd3695:data <=32'hFFFEFFAB;
14'd3696:data <=32'hFFF5FF9C;14'd3697:data <=32'hFFE4FF8F;14'd3698:data <=32'hFFCFFF87;
14'd3699:data <=32'hFFB5FF88;14'd3700:data <=32'hFF9CFF90;14'd3701:data <=32'hFF89FF9E;
14'd3702:data <=32'hFF78FFB0;14'd3703:data <=32'hFF6DFFC3;14'd3704:data <=32'hFF65FFD6;
14'd3705:data <=32'hFF60FFE8;14'd3706:data <=32'hFF5CFFFB;14'd3707:data <=32'hFF59000E;
14'd3708:data <=32'hFF590023;14'd3709:data <=32'hFF5D0038;14'd3710:data <=32'hFF64004D;
14'd3711:data <=32'hFF6F005E;14'd3712:data <=32'hFF3E00BF;14'd3713:data <=32'hFF5F00E8;
14'd3714:data <=32'hFF8300EE;14'd3715:data <=32'hFF6A0070;14'd3716:data <=32'hFF500052;
14'd3717:data <=32'hFF4D0077;14'd3718:data <=32'hFF5600A0;14'd3719:data <=32'hFF6B00CB;
14'd3720:data <=32'hFF9000F1;14'd3721:data <=32'hFFC0010C;14'd3722:data <=32'hFFF80118;
14'd3723:data <=32'h00310116;14'd3724:data <=32'h00670105;14'd3725:data <=32'h009400E8;
14'd3726:data <=32'h00BA00C2;14'd3727:data <=32'h00D50096;14'd3728:data <=32'h00E50067;
14'd3729:data <=32'h00EC0036;14'd3730:data <=32'h00E60005;14'd3731:data <=32'h00D5FFD6;
14'd3732:data <=32'h00B8FFB0;14'd3733:data <=32'h0091FF94;14'd3734:data <=32'h0067FF85;
14'd3735:data <=32'h003CFF86;14'd3736:data <=32'h0018FF92;14'd3737:data <=32'hFFFDFFA8;
14'd3738:data <=32'hFFEEFFC3;14'd3739:data <=32'hFFE9FFDC;14'd3740:data <=32'hFFEDFFF2;
14'd3741:data <=32'hFFF40003;14'd3742:data <=32'h0000000D;14'd3743:data <=32'h000A0014;
14'd3744:data <=32'h00150019;14'd3745:data <=32'h0021001B;14'd3746:data <=32'h002D001C;
14'd3747:data <=32'h003B001A;14'd3748:data <=32'h00480013;14'd3749:data <=32'h0055000A;
14'd3750:data <=32'h005EFFFC;14'd3751:data <=32'h0065FFEB;14'd3752:data <=32'h0067FFDA;
14'd3753:data <=32'h0066FFC8;14'd3754:data <=32'h0061FFB8;14'd3755:data <=32'h005CFFA8;
14'd3756:data <=32'h0055FF99;14'd3757:data <=32'h004CFF8A;14'd3758:data <=32'h003EFF79;
14'd3759:data <=32'h002CFF68;14'd3760:data <=32'h0015FF5B;14'd3761:data <=32'hFFF8FF54;
14'd3762:data <=32'hFFD8FF54;14'd3763:data <=32'hFFB8FF5E;14'd3764:data <=32'hFF9DFF72;
14'd3765:data <=32'hFF8AFF8C;14'd3766:data <=32'hFF80FFA7;14'd3767:data <=32'hFF80FFC1;
14'd3768:data <=32'hFF88FFD8;14'd3769:data <=32'hFF93FFE6;14'd3770:data <=32'hFF9FFFEE;
14'd3771:data <=32'hFFA8FFF0;14'd3772:data <=32'hFFAFFFEE;14'd3773:data <=32'hFFB2FFEB;
14'd3774:data <=32'hFFB1FFE5;14'd3775:data <=32'hFFADFFDF;14'd3776:data <=32'hFF2EFFE7;
14'd3777:data <=32'hFF200009;14'd3778:data <=32'hFF310028;14'd3779:data <=32'hFF96FFF4;
14'd3780:data <=32'hFF69FFC2;14'd3781:data <=32'hFF4CFFD7;14'd3782:data <=32'hFF34FFF8;
14'd3783:data <=32'hFF250022;14'd3784:data <=32'hFF230052;14'd3785:data <=32'hFF330082;
14'd3786:data <=32'hFF4E00AB;14'd3787:data <=32'hFF7300C9;14'd3788:data <=32'hFF9C00DE;
14'd3789:data <=32'hFFC700E7;14'd3790:data <=32'hFFF100E8;14'd3791:data <=32'h001800E1;
14'd3792:data <=32'h003E00D3;14'd3793:data <=32'h005D00BE;14'd3794:data <=32'h007A00A3;
14'd3795:data <=32'h008E0083;14'd3796:data <=32'h0098005F;14'd3797:data <=32'h0099003C;
14'd3798:data <=32'h0091001C;14'd3799:data <=32'h00810004;14'd3800:data <=32'h006FFFF3;
14'd3801:data <=32'h005DFFEA;14'd3802:data <=32'h004EFFE5;14'd3803:data <=32'h0041FFE3;
14'd3804:data <=32'h0037FFE2;14'd3805:data <=32'h002DFFDF;14'd3806:data <=32'h0022FFDF;
14'd3807:data <=32'h0015FFE0;14'd3808:data <=32'h0007FFE6;14'd3809:data <=32'hFFF9FFF1;
14'd3810:data <=32'hFFF10002;14'd3811:data <=32'hFFEF0016;14'd3812:data <=32'hFFF4002C;
14'd3813:data <=32'h0002003E;14'd3814:data <=32'h0016004C;14'd3815:data <=32'h002E0053;
14'd3816:data <=32'h00480055;14'd3817:data <=32'h0063004F;14'd3818:data <=32'h007C0042;
14'd3819:data <=32'h0093002E;14'd3820:data <=32'h00A80014;14'd3821:data <=32'h00B7FFF4;
14'd3822:data <=32'h00BFFFCF;14'd3823:data <=32'h00BCFFA5;14'd3824:data <=32'h00AFFF7B;
14'd3825:data <=32'h0093FF55;14'd3826:data <=32'h006EFF38;14'd3827:data <=32'h0042FF26;
14'd3828:data <=32'h0013FF24;14'd3829:data <=32'hFFE8FF2D;14'd3830:data <=32'hFFC5FF42;
14'd3831:data <=32'hFFAEFF5C;14'd3832:data <=32'hFF9FFF78;14'd3833:data <=32'hFF9AFF92;
14'd3834:data <=32'hFF9CFFA7;14'd3835:data <=32'hFFA0FFB7;14'd3836:data <=32'hFFA5FFC2;
14'd3837:data <=32'hFFABFFC8;14'd3838:data <=32'hFFB1FFCD;14'd3839:data <=32'hFFB5FFCC;
14'd3840:data <=32'hFFC7FFB2;14'd3841:data <=32'hFFB9FFA6;14'd3842:data <=32'hFFA6FFAE;
14'd3843:data <=32'hFF93FFE3;14'd3844:data <=32'hFF77FFB0;14'd3845:data <=32'hFF66FFBE;
14'd3846:data <=32'hFF56FFD3;14'd3847:data <=32'hFF4BFFEE;14'd3848:data <=32'hFF47000E;
14'd3849:data <=32'hFF50002E;14'd3850:data <=32'hFF5F004A;14'd3851:data <=32'hFF74005D;
14'd3852:data <=32'hFF8C0069;14'd3853:data <=32'hFFA2006F;14'd3854:data <=32'hFFB30070;
14'd3855:data <=32'hFFC0006F;14'd3856:data <=32'hFFCC006E;14'd3857:data <=32'hFFD6006E;
14'd3858:data <=32'hFFE1006E;14'd3859:data <=32'hFFEC006D;14'd3860:data <=32'hFFF6006B;
14'd3861:data <=32'hFFFF0067;14'd3862:data <=32'h00060064;14'd3863:data <=32'h000B0062;
14'd3864:data <=32'h00130062;14'd3865:data <=32'h001B0063;14'd3866:data <=32'h00280061;
14'd3867:data <=32'h0037005D;14'd3868:data <=32'h00470053;14'd3869:data <=32'h00530042;
14'd3870:data <=32'h005B002B;14'd3871:data <=32'h005A0013;14'd3872:data <=32'h004EFFFD;
14'd3873:data <=32'h003CFFED;14'd3874:data <=32'h0025FFE4;14'd3875:data <=32'h000EFFE7;
14'd3876:data <=32'hFFFAFFF2;14'd3877:data <=32'hFFEC0003;14'd3878:data <=32'hFFE40018;
14'd3879:data <=32'hFFE5002F;14'd3880:data <=32'hFFED0044;14'd3881:data <=32'hFFFB0058;
14'd3882:data <=32'h000E0069;14'd3883:data <=32'h00270073;14'd3884:data <=32'h00440078;
14'd3885:data <=32'h00640074;14'd3886:data <=32'h00860068;14'd3887:data <=32'h00A30051;
14'd3888:data <=32'h00BB0032;14'd3889:data <=32'h00C7000D;14'd3890:data <=32'h00CAFFE5;
14'd3891:data <=32'h00C2FFC0;14'd3892:data <=32'h00B1FFA1;14'd3893:data <=32'h009AFF89;
14'd3894:data <=32'h0084FF79;14'd3895:data <=32'h0070FF6F;14'd3896:data <=32'h005DFF67;
14'd3897:data <=32'h004DFF5F;14'd3898:data <=32'h003EFF57;14'd3899:data <=32'h002BFF4E;
14'd3900:data <=32'h0017FF46;14'd3901:data <=32'hFFFFFF42;14'd3902:data <=32'hFFE6FF42;
14'd3903:data <=32'hFFCDFF45;14'd3904:data <=32'hFFE1FFDF;14'd3905:data <=32'hFFF2FFD2;
14'd3906:data <=32'hFFF2FFB5;14'd3907:data <=32'hFF94FF55;14'd3908:data <=32'hFF65FF31;
14'd3909:data <=32'hFF42FF50;14'd3910:data <=32'hFF27FF78;14'd3911:data <=32'hFF16FFA7;
14'd3912:data <=32'hFF12FFD9;14'd3913:data <=32'hFF1D000B;14'd3914:data <=32'hFF350036;
14'd3915:data <=32'hFF570054;14'd3916:data <=32'hFF7D0065;14'd3917:data <=32'hFFA20068;
14'd3918:data <=32'hFFC0005F;14'd3919:data <=32'hFFD50052;14'd3920:data <=32'hFFE20041;
14'd3921:data <=32'hFFE90032;14'd3922:data <=32'hFFE80025;14'd3923:data <=32'hFFE4001A;
14'd3924:data <=32'hFFDD0013;14'd3925:data <=32'hFFD30010;14'd3926:data <=32'hFFC90011;
14'd3927:data <=32'hFFBD0017;14'd3928:data <=32'hFFB40024;14'd3929:data <=32'hFFB00035;
14'd3930:data <=32'hFFB3004A;14'd3931:data <=32'hFFBF005D;14'd3932:data <=32'hFFD2006C;
14'd3933:data <=32'hFFEA0072;14'd3934:data <=32'h0002006F;14'd3935:data <=32'h00150065;
14'd3936:data <=32'h00240055;14'd3937:data <=32'h002A0044;14'd3938:data <=32'h00290033;
14'd3939:data <=32'h00230027;14'd3940:data <=32'h001B0020;14'd3941:data <=32'h0012001E;
14'd3942:data <=32'h000C001F;14'd3943:data <=32'h00070021;14'd3944:data <=32'h00030026;
14'd3945:data <=32'h0000002C;14'd3946:data <=32'hFFFF0033;14'd3947:data <=32'hFFFF003B;
14'd3948:data <=32'h00020045;14'd3949:data <=32'h00080050;14'd3950:data <=32'h00130058;
14'd3951:data <=32'h00220060;14'd3952:data <=32'h00310062;14'd3953:data <=32'h00420060;
14'd3954:data <=32'h0051005C;14'd3955:data <=32'h005E0056;14'd3956:data <=32'h006A004F;
14'd3957:data <=32'h0076004A;14'd3958:data <=32'h00850046;14'd3959:data <=32'h0098003F;
14'd3960:data <=32'h00AE0032;14'd3961:data <=32'h00C7001D;14'd3962:data <=32'h00DDFFFD;
14'd3963:data <=32'h00EBFFD6;14'd3964:data <=32'h00EEFFA6;14'd3965:data <=32'h00E5FF74;
14'd3966:data <=32'h00CFFF45;14'd3967:data <=32'h00AEFF1B;14'd3968:data <=32'h000CFFA4;
14'd3969:data <=32'h0016FF9F;14'd3970:data <=32'h0031FF8D;14'd3971:data <=32'h006CFF0E;
14'd3972:data <=32'h002AFEC3;14'd3973:data <=32'hFFEAFEC3;14'd3974:data <=32'hFFABFED4;
14'd3975:data <=32'hFF74FEF3;14'd3976:data <=32'hFF47FF20;14'd3977:data <=32'hFF29FF56;
14'd3978:data <=32'hFF1EFF91;14'd3979:data <=32'hFF23FFC6;14'd3980:data <=32'hFF35FFF2;
14'd3981:data <=32'hFF500013;14'd3982:data <=32'hFF6D0027;14'd3983:data <=32'hFF880032;
14'd3984:data <=32'hFF9F0035;14'd3985:data <=32'hFFB30034;14'd3986:data <=32'hFFC20030;
14'd3987:data <=32'hFFCF002A;14'd3988:data <=32'hFFD90022;14'd3989:data <=32'hFFDF0018;
14'd3990:data <=32'hFFE0000E;14'd3991:data <=32'hFFDC0005;14'd3992:data <=32'hFFD40001;
14'd3993:data <=32'hFFCC0000;14'd3994:data <=32'hFFC30005;14'd3995:data <=32'hFFBF000D;
14'd3996:data <=32'hFFBE0017;14'd3997:data <=32'hFFC20020;14'd3998:data <=32'hFFC80024;
14'd3999:data <=32'hFFCD0026;14'd4000:data <=32'hFFCF0026;14'd4001:data <=32'hFFCF0025;
14'd4002:data <=32'hFFCC0027;14'd4003:data <=32'hFFC8002D;14'd4004:data <=32'hFFC60036;
14'd4005:data <=32'hFFC70042;14'd4006:data <=32'hFFCE004E;14'd4007:data <=32'hFFD90057;
14'd4008:data <=32'hFFE7005E;14'd4009:data <=32'hFFF6005E;14'd4010:data <=32'h0003005B;
14'd4011:data <=32'h000D0055;14'd4012:data <=32'h0013004D;14'd4013:data <=32'h00170045;
14'd4014:data <=32'h0018003E;14'd4015:data <=32'h00170038;14'd4016:data <=32'h00130034;
14'd4017:data <=32'h00100033;14'd4018:data <=32'h00080033;14'd4019:data <=32'h00010039;
14'd4020:data <=32'hFFFB0045;14'd4021:data <=32'hFFF70057;14'd4022:data <=32'hFFFC006E;
14'd4023:data <=32'h000C0088;14'd4024:data <=32'h0028009E;14'd4025:data <=32'h004F00AD;
14'd4026:data <=32'h007E00AE;14'd4027:data <=32'h00AF00A0;14'd4028:data <=32'h00DB0082;
14'd4029:data <=32'h01000058;14'd4030:data <=32'h01170025;14'd4031:data <=32'h0123FFEE;
14'd4032:data <=32'h00A9FFEA;14'd4033:data <=32'h00BFFFD0;14'd4034:data <=32'h00D0FFC2;
14'd4035:data <=32'h00FAFFCB;14'd4036:data <=32'h00DDFF64;14'd4037:data <=32'h00BBFF3F;
14'd4038:data <=32'h0092FF25;14'd4039:data <=32'h0065FF15;14'd4040:data <=32'h0036FF10;
14'd4041:data <=32'h000BFF19;14'd4042:data <=32'hFFE8FF2B;14'd4043:data <=32'hFFCEFF40;
14'd4044:data <=32'hFFBDFF56;14'd4045:data <=32'hFFB2FF69;14'd4046:data <=32'hFFA9FF78;
14'd4047:data <=32'hFF9FFF86;14'd4048:data <=32'hFF95FF92;14'd4049:data <=32'hFF8BFFA2;
14'd4050:data <=32'hFF82FFB6;14'd4051:data <=32'hFF7EFFCC;14'd4052:data <=32'hFF7FFFE2;
14'd4053:data <=32'hFF86FFF7;14'd4054:data <=32'hFF900008;14'd4055:data <=32'hFF9D0014;
14'd4056:data <=32'hFFAA001E;14'd4057:data <=32'hFFB80024;14'd4058:data <=32'hFFC60027;
14'd4059:data <=32'hFFD40029;14'd4060:data <=32'hFFE30026;14'd4061:data <=32'hFFF0001F;
14'd4062:data <=32'hFFFD0012;14'd4063:data <=32'h00020001;14'd4064:data <=32'h0000FFEE;
14'd4065:data <=32'hFFF6FFDB;14'd4066:data <=32'hFFE3FFCE;14'd4067:data <=32'hFFCBFFC9;
14'd4068:data <=32'hFFB2FFCE;14'd4069:data <=32'hFF9CFFDD;14'd4070:data <=32'hFF8DFFF1;
14'd4071:data <=32'hFF85000B;14'd4072:data <=32'hFF870024;14'd4073:data <=32'hFF8F003C;
14'd4074:data <=32'hFF9B004D;14'd4075:data <=32'hFFAB0059;14'd4076:data <=32'hFFBC0061;
14'd4077:data <=32'hFFCB0067;14'd4078:data <=32'hFFDB0067;14'd4079:data <=32'hFFE80065;
14'd4080:data <=32'hFFF3005F;14'd4081:data <=32'hFFFA0059;14'd4082:data <=32'hFFFE0050;
14'd4083:data <=32'hFFFD004A;14'd4084:data <=32'hFFF70047;14'd4085:data <=32'hFFEF004B;
14'd4086:data <=32'hFFE70056;14'd4087:data <=32'hFFE60069;14'd4088:data <=32'hFFED007F;
14'd4089:data <=32'hFFFF0095;14'd4090:data <=32'h001A00A6;14'd4091:data <=32'h003C00AD;
14'd4092:data <=32'h006100AA;14'd4093:data <=32'h0083009C;14'd4094:data <=32'h00A10086;
14'd4095:data <=32'h00B7006B;14'd4096:data <=32'h008300BD;14'd4097:data <=32'h00C100B3;
14'd4098:data <=32'h00E50098;14'd4099:data <=32'h00A10050;14'd4100:data <=32'h009C0002;
14'd4101:data <=32'h0098FFF2;14'd4102:data <=32'h0092FFE3;14'd4103:data <=32'h008BFFD6;
14'd4104:data <=32'h0083FFCC;14'd4105:data <=32'h007CFFC6;14'd4106:data <=32'h0078FFC0;
14'd4107:data <=32'h0077FFB9;14'd4108:data <=32'h0079FFAE;14'd4109:data <=32'h007BFF9D;
14'd4110:data <=32'h0076FF85;14'd4111:data <=32'h006BFF6B;14'd4112:data <=32'h0054FF52;
14'd4113:data <=32'h0034FF3E;14'd4114:data <=32'h000EFF35;14'd4115:data <=32'hFFE6FF37;
14'd4116:data <=32'hFFC0FF45;14'd4117:data <=32'hFFA1FF5B;14'd4118:data <=32'hFF89FF77;
14'd4119:data <=32'hFF7AFF96;14'd4120:data <=32'hFF72FFB6;14'd4121:data <=32'hFF71FFD7;
14'd4122:data <=32'hFF79FFF6;14'd4123:data <=32'hFF880012;14'd4124:data <=32'hFF9D0028;
14'd4125:data <=32'hFFB90038;14'd4126:data <=32'hFFD8003C;14'd4127:data <=32'hFFF60035;
14'd4128:data <=32'h000F0025;14'd4129:data <=32'h001F000C;14'd4130:data <=32'h0023FFF0;
14'd4131:data <=32'h001EFFD5;14'd4132:data <=32'h000FFFBF;14'd4133:data <=32'hFFFAFFB1;
14'd4134:data <=32'hFFE3FFAB;14'd4135:data <=32'hFFCDFFAC;14'd4136:data <=32'hFFBAFFB3;
14'd4137:data <=32'hFFABFFBC;14'd4138:data <=32'hFF9EFFC5;14'd4139:data <=32'hFF92FFD1;
14'd4140:data <=32'hFF87FFDE;14'd4141:data <=32'hFF7EFFEC;14'd4142:data <=32'hFF76FFFE;
14'd4143:data <=32'hFF700011;14'd4144:data <=32'hFF700026;14'd4145:data <=32'hFF73003C;
14'd4146:data <=32'hFF78004D;14'd4147:data <=32'hFF800060;14'd4148:data <=32'hFF8A0070;
14'd4149:data <=32'hFF940081;14'd4150:data <=32'hFFA00093;14'd4151:data <=32'hFFB000A6;
14'd4152:data <=32'hFFC500B7;14'd4153:data <=32'hFFE300C7;14'd4154:data <=32'h000500CF;
14'd4155:data <=32'h002B00CE;14'd4156:data <=32'h005000C2;14'd4157:data <=32'h007000AB;
14'd4158:data <=32'h0087008D;14'd4159:data <=32'h0092006E;14'd4160:data <=32'hFFCF00CA;
14'd4161:data <=32'h000000F1;14'd4162:data <=32'h004100F4;14'd4163:data <=32'h00810059;
14'd4164:data <=32'h0072000D;14'd4165:data <=32'h00610006;14'd4166:data <=32'h00520004;
14'd4167:data <=32'h00460007;14'd4168:data <=32'h003E000E;14'd4169:data <=32'h003B0019;
14'd4170:data <=32'h00400027;14'd4171:data <=32'h004D0033;14'd4172:data <=32'h00630038;
14'd4173:data <=32'h007E0031;14'd4174:data <=32'h00970020;14'd4175:data <=32'h00AC0003;
14'd4176:data <=32'h00B4FFDD;14'd4177:data <=32'h00B2FFB6;14'd4178:data <=32'h00A2FF91;
14'd4179:data <=32'h0088FF74;14'd4180:data <=32'h0069FF5E;14'd4181:data <=32'h0047FF53;
14'd4182:data <=32'h0026FF50;14'd4183:data <=32'h0005FF54;14'd4184:data <=32'hFFE8FF5E;
14'd4185:data <=32'hFFCDFF6D;14'd4186:data <=32'hFFB9FF82;14'd4187:data <=32'hFFA8FF9B;
14'd4188:data <=32'hFFA0FFB7;14'd4189:data <=32'hFFA0FFD3;14'd4190:data <=32'hFFAAFFEC;
14'd4191:data <=32'hFFB90000;14'd4192:data <=32'hFFCD000B;14'd4193:data <=32'hFFE1000F;
14'd4194:data <=32'hFFF3000C;14'd4195:data <=32'h00000004;14'd4196:data <=32'h0008FFFB;
14'd4197:data <=32'h000EFFF1;14'd4198:data <=32'h0010FFE8;14'd4199:data <=32'h0014FFE0;
14'd4200:data <=32'h0017FFD6;14'd4201:data <=32'h0019FFC8;14'd4202:data <=32'h0017FFB8;
14'd4203:data <=32'h0011FFA4;14'd4204:data <=32'h0004FF90;14'd4205:data <=32'hFFEFFF7E;
14'd4206:data <=32'hFFD1FF71;14'd4207:data <=32'hFFB0FF6D;14'd4208:data <=32'hFF8BFF72;
14'd4209:data <=32'hFF68FF7F;14'd4210:data <=32'hFF48FF97;14'd4211:data <=32'hFF2DFFB4;
14'd4212:data <=32'hFF17FFD9;14'd4213:data <=32'hFF080003;14'd4214:data <=32'hFF010032;
14'd4215:data <=32'hFF050065;14'd4216:data <=32'hFF150097;14'd4217:data <=32'hFF3400C8;
14'd4218:data <=32'hFF5F00F0;14'd4219:data <=32'hFF96010A;14'd4220:data <=32'hFFD00115;
14'd4221:data <=32'h000A010E;14'd4222:data <=32'h003D00F8;14'd4223:data <=32'h006300D6;
14'd4224:data <=32'hFFB5007B;14'd4225:data <=32'hFFC1009F;14'd4226:data <=32'hFFE300C6;
14'd4227:data <=32'h005E00CA;14'd4228:data <=32'h00670075;14'd4229:data <=32'h00660060;
14'd4230:data <=32'h0063004E;14'd4231:data <=32'h005E0040;14'd4232:data <=32'h00560037;
14'd4233:data <=32'h004E0033;14'd4234:data <=32'h00480034;14'd4235:data <=32'h00480039;
14'd4236:data <=32'h004E003F;14'd4237:data <=32'h005A0041;14'd4238:data <=32'h006B003C;
14'd4239:data <=32'h007B0030;14'd4240:data <=32'h0086001C;14'd4241:data <=32'h008B0005;
14'd4242:data <=32'h0088FFED;14'd4243:data <=32'h007EFFDA;14'd4244:data <=32'h0071FFCB;
14'd4245:data <=32'h0064FFC1;14'd4246:data <=32'h0056FFBC;14'd4247:data <=32'h004CFFB8;
14'd4248:data <=32'h0042FFB5;14'd4249:data <=32'h003AFFB2;14'd4250:data <=32'h0030FFAF;
14'd4251:data <=32'h0025FFAE;14'd4252:data <=32'h001BFFAE;14'd4253:data <=32'h0011FFB2;
14'd4254:data <=32'h0009FFB7;14'd4255:data <=32'h0005FFBC;14'd4256:data <=32'h0000FFC1;
14'd4257:data <=32'hFFFEFFC4;14'd4258:data <=32'hFFF9FFC5;14'd4259:data <=32'hFFF5FFCA;
14'd4260:data <=32'hFFEEFFCE;14'd4261:data <=32'hFFE9FFD7;14'd4262:data <=32'hFFE8FFE4;
14'd4263:data <=32'hFFEEFFF1;14'd4264:data <=32'hFFF9FFFC;14'd4265:data <=32'h000C0002;
14'd4266:data <=32'h0021FFFF;14'd4267:data <=32'h0036FFF3;14'd4268:data <=32'h0046FFDC;
14'd4269:data <=32'h004FFFBF;14'd4270:data <=32'h004DFF9D;14'd4271:data <=32'h003FFF7D;
14'd4272:data <=32'h0028FF60;14'd4273:data <=32'h0008FF4A;14'd4274:data <=32'hFFE2FF3C;
14'd4275:data <=32'hFFB9FF35;14'd4276:data <=32'hFF8CFF3A;14'd4277:data <=32'hFF60FF49;
14'd4278:data <=32'hFF35FF62;14'd4279:data <=32'hFF11FF87;14'd4280:data <=32'hFEF5FFB7;
14'd4281:data <=32'hFEE5FFEE;14'd4282:data <=32'hFEE60027;14'd4283:data <=32'hFEF6005E;
14'd4284:data <=32'hFF14008D;14'd4285:data <=32'hFF3A00B0;14'd4286:data <=32'hFF6500C6;
14'd4287:data <=32'hFF8F00CF;14'd4288:data <=32'hFF91009A;14'd4289:data <=32'hFFA000B0;
14'd4290:data <=32'hFFA600C7;14'd4291:data <=32'hFF8300DD;14'd4292:data <=32'hFF9C00AE;
14'd4293:data <=32'hFFB300BB;14'd4294:data <=32'hFFCD00C4;14'd4295:data <=32'hFFE900CA;
14'd4296:data <=32'h000500CA;14'd4297:data <=32'h002100C4;14'd4298:data <=32'h003A00BD;
14'd4299:data <=32'h005200B1;14'd4300:data <=32'h006900A4;14'd4301:data <=32'h00810090;
14'd4302:data <=32'h00960077;14'd4303:data <=32'h00A60059;14'd4304:data <=32'h00AD0035;
14'd4305:data <=32'h00AA0010;14'd4306:data <=32'h009BFFEE;14'd4307:data <=32'h0083FFD4;
14'd4308:data <=32'h0067FFC5;14'd4309:data <=32'h004AFFC2;14'd4310:data <=32'h0032FFC8;
14'd4311:data <=32'h001FFFD4;14'd4312:data <=32'h0017FFE2;14'd4313:data <=32'h0013FFF1;
14'd4314:data <=32'h0016FFFD;14'd4315:data <=32'h001B0005;14'd4316:data <=32'h0024000B;
14'd4317:data <=32'h002C000D;14'd4318:data <=32'h0036000D;14'd4319:data <=32'h00400008;
14'd4320:data <=32'h0049FFFF;14'd4321:data <=32'h0050FFF3;14'd4322:data <=32'h0052FFE4;
14'd4323:data <=32'h004DFFD4;14'd4324:data <=32'h0044FFC6;14'd4325:data <=32'h0035FFBF;
14'd4326:data <=32'h0026FFBE;14'd4327:data <=32'h0018FFC3;14'd4328:data <=32'h000FFFCD;
14'd4329:data <=32'h0010FFDA;14'd4330:data <=32'h0016FFE4;14'd4331:data <=32'h0022FFE8;
14'd4332:data <=32'h002FFFE5;14'd4333:data <=32'h003CFFDB;14'd4334:data <=32'h0045FFCC;
14'd4335:data <=32'h0047FFB9;14'd4336:data <=32'h0044FFA6;14'd4337:data <=32'h003CFF93;
14'd4338:data <=32'h002FFF81;14'd4339:data <=32'h001FFF73;14'd4340:data <=32'h000BFF66;
14'd4341:data <=32'hFFF4FF5D;14'd4342:data <=32'hFFDAFF58;14'd4343:data <=32'hFFBDFF58;
14'd4344:data <=32'hFFA0FF60;14'd4345:data <=32'hFF85FF6E;14'd4346:data <=32'hFF6EFF83;
14'd4347:data <=32'hFF5EFF9B;14'd4348:data <=32'hFF56FFB3;14'd4349:data <=32'hFF52FFCA;
14'd4350:data <=32'hFF50FFDB;14'd4351:data <=32'hFF4EFFEB;14'd4352:data <=32'hFF130038;
14'd4353:data <=32'hFF16005F;14'd4354:data <=32'hFF24006F;14'd4355:data <=32'hFF23FFFD;
14'd4356:data <=32'hFF13FFE5;14'd4357:data <=32'hFF05000F;14'd4358:data <=32'hFF020040;
14'd4359:data <=32'hFF0B0072;14'd4360:data <=32'hFF2100A0;14'd4361:data <=32'hFF3F00C7;
14'd4362:data <=32'hFF6600E8;14'd4363:data <=32'hFF930101;14'd4364:data <=32'hFFC60110;
14'd4365:data <=32'hFFFC0115;14'd4366:data <=32'h0033010A;14'd4367:data <=32'h006600F3;
14'd4368:data <=32'h009200CD;14'd4369:data <=32'h00B0009C;14'd4370:data <=32'h00BE0068;
14'd4371:data <=32'h00BA0034;14'd4372:data <=32'h00A90009;14'd4373:data <=32'h008FFFE9;
14'd4374:data <=32'h006FFFD5;14'd4375:data <=32'h0050FFCD;14'd4376:data <=32'h0034FFCD;
14'd4377:data <=32'h001FFFD5;14'd4378:data <=32'h000EFFDF;14'd4379:data <=32'h0002FFEC;
14'd4380:data <=32'hFFFAFFFB;14'd4381:data <=32'hFFF7000B;14'd4382:data <=32'hFFF8001B;
14'd4383:data <=32'hFFFF0029;14'd4384:data <=32'h000C0035;14'd4385:data <=32'h001B003C;
14'd4386:data <=32'h002C003E;14'd4387:data <=32'h003B0039;14'd4388:data <=32'h00480030;
14'd4389:data <=32'h00510027;14'd4390:data <=32'h0055001D;14'd4391:data <=32'h00590014;
14'd4392:data <=32'h005D000E;14'd4393:data <=32'h00620008;14'd4394:data <=32'h00690000;
14'd4395:data <=32'h0072FFF5;14'd4396:data <=32'h0079FFE5;14'd4397:data <=32'h007DFFD0;
14'd4398:data <=32'h007AFFBA;14'd4399:data <=32'h006FFFA3;14'd4400:data <=32'h0060FF90;
14'd4401:data <=32'h004CFF83;14'd4402:data <=32'h0034FF7B;14'd4403:data <=32'h0021FF7A;
14'd4404:data <=32'h000EFF7E;14'd4405:data <=32'h0000FF84;14'd4406:data <=32'hFFF4FF8B;
14'd4407:data <=32'hFFEBFF92;14'd4408:data <=32'hFFE4FF9A;14'd4409:data <=32'hFFE0FFA1;
14'd4410:data <=32'hFFDFFFA8;14'd4411:data <=32'hFFE1FFAC;14'd4412:data <=32'hFFE5FFAD;
14'd4413:data <=32'hFFEAFFA6;14'd4414:data <=32'hFFECFF9A;14'd4415:data <=32'hFFE5FF88;
14'd4416:data <=32'hFF65FF75;14'd4417:data <=32'hFF47FF83;14'd4418:data <=32'hFF42FF9C;
14'd4419:data <=32'hFFA9FF83;14'd4420:data <=32'hFF89FF4A;14'd4421:data <=32'hFF5DFF59;
14'd4422:data <=32'hFF35FF75;14'd4423:data <=32'hFF17FF9D;14'd4424:data <=32'hFF04FFC9;
14'd4425:data <=32'hFEFAFFF8;14'd4426:data <=32'hFEFB0029;14'd4427:data <=32'hFF050058;
14'd4428:data <=32'hFF1B0085;14'd4429:data <=32'hFF3A00AE;14'd4430:data <=32'hFF6400CD;
14'd4431:data <=32'hFF9300E2;14'd4432:data <=32'hFFC600E7;14'd4433:data <=32'hFFF700DE;
14'd4434:data <=32'h002000CA;14'd4435:data <=32'h003D00AE;14'd4436:data <=32'h0050008F;
14'd4437:data <=32'h00590072;14'd4438:data <=32'h005B0058;14'd4439:data <=32'h00580043;
14'd4440:data <=32'h00550032;14'd4441:data <=32'h00500024;14'd4442:data <=32'h004B0015;
14'd4443:data <=32'h00410008;14'd4444:data <=32'h0036FFFC;14'd4445:data <=32'h0027FFF5;
14'd4446:data <=32'h0018FFF1;14'd4447:data <=32'h0007FFF5;14'd4448:data <=32'hFFFAFFFC;
14'd4449:data <=32'hFFEF0008;14'd4450:data <=32'hFFE90016;14'd4451:data <=32'hFFE70024;
14'd4452:data <=32'hFFE80034;14'd4453:data <=32'hFFEC0042;14'd4454:data <=32'hFFF40052;
14'd4455:data <=32'h00000062;14'd4456:data <=32'h00110071;14'd4457:data <=32'h002A007B;
14'd4458:data <=32'h00490081;14'd4459:data <=32'h006A007C;14'd4460:data <=32'h008D006E;
14'd4461:data <=32'h00AB0054;14'd4462:data <=32'h00C20031;14'd4463:data <=32'h00CC0007;
14'd4464:data <=32'h00CAFFDD;14'd4465:data <=32'h00BDFFB6;14'd4466:data <=32'h00A7FF96;
14'd4467:data <=32'h008BFF80;14'd4468:data <=32'h006DFF72;14'd4469:data <=32'h0050FF6D;
14'd4470:data <=32'h0036FF6D;14'd4471:data <=32'h001EFF73;14'd4472:data <=32'h000CFF7D;
14'd4473:data <=32'hFFFDFF8B;14'd4474:data <=32'hFFF5FF9A;14'd4475:data <=32'hFFF3FFA9;
14'd4476:data <=32'hFFF8FFB5;14'd4477:data <=32'h0004FFBA;14'd4478:data <=32'h0011FFB7;
14'd4479:data <=32'h001CFFA9;14'd4480:data <=32'h0022FF91;14'd4481:data <=32'h001AFF73;
14'd4482:data <=32'h0003FF69;14'd4483:data <=32'hFFE3FF93;14'd4484:data <=32'hFFD4FF53;
14'd4485:data <=32'hFFB6FF58;14'd4486:data <=32'hFF99FF64;14'd4487:data <=32'hFF81FF78;
14'd4488:data <=32'hFF70FF8F;14'd4489:data <=32'hFF64FFA7;14'd4490:data <=32'hFF5CFFBE;
14'd4491:data <=32'hFF58FFD5;14'd4492:data <=32'hFF56FFED;14'd4493:data <=32'hFF590005;
14'd4494:data <=32'hFF60001D;14'd4495:data <=32'hFF6D0031;14'd4496:data <=32'hFF7D0041;
14'd4497:data <=32'hFF8E004B;14'd4498:data <=32'hFF9E0050;14'd4499:data <=32'hFFAA0051;
14'd4500:data <=32'hFFB30051;14'd4501:data <=32'hFFB80054;14'd4502:data <=32'hFFBC005B;
14'd4503:data <=32'hFFC40064;14'd4504:data <=32'hFFD0006E;14'd4505:data <=32'hFFE20076;
14'd4506:data <=32'hFFF80078;14'd4507:data <=32'h000F0072;14'd4508:data <=32'h00230065;
14'd4509:data <=32'h00310053;14'd4510:data <=32'h0039003D;14'd4511:data <=32'h00390028;
14'd4512:data <=32'h00320015;14'd4513:data <=32'h00270006;14'd4514:data <=32'h0018FFFB;
14'd4515:data <=32'h0007FFF5;14'd4516:data <=32'hFFF4FFF4;14'd4517:data <=32'hFFE1FFFA;
14'd4518:data <=32'hFFCE0007;14'd4519:data <=32'hFFC0001B;14'd4520:data <=32'hFFB60036;
14'd4521:data <=32'hFFB70054;14'd4522:data <=32'hFFC30074;14'd4523:data <=32'hFFDA0091;
14'd4524:data <=32'hFFFB00A5;14'd4525:data <=32'h002200AF;14'd4526:data <=32'h004900AB;
14'd4527:data <=32'h006F009D;14'd4528:data <=32'h008C0086;14'd4529:data <=32'h00A1006A;
14'd4530:data <=32'h00AF004C;14'd4531:data <=32'h00B6002F;14'd4532:data <=32'h00B70015;
14'd4533:data <=32'h00B5FFFD;14'd4534:data <=32'h00B1FFE6;14'd4535:data <=32'h00AAFFD1;
14'd4536:data <=32'h00A0FFBD;14'd4537:data <=32'h0095FFAC;14'd4538:data <=32'h0087FF9C;
14'd4539:data <=32'h0079FF92;14'd4540:data <=32'h006CFF8A;14'd4541:data <=32'h0062FF83;
14'd4542:data <=32'h0059FF7A;14'd4543:data <=32'h0051FF6E;14'd4544:data <=32'h002AFFF9;
14'd4545:data <=32'h004BFFE8;14'd4546:data <=32'h0058FFC1;14'd4547:data <=32'h0017FF47;
14'd4548:data <=32'hFFF9FF0B;14'd4549:data <=32'hFFCAFF18;14'd4550:data <=32'hFFA3FF30;
14'd4551:data <=32'hFF84FF52;14'd4552:data <=32'hFF73FF77;14'd4553:data <=32'hFF6DFF9C;
14'd4554:data <=32'hFF71FFBB;14'd4555:data <=32'hFF7AFFD5;14'd4556:data <=32'hFF87FFE9;
14'd4557:data <=32'hFF96FFF8;14'd4558:data <=32'hFFA50001;14'd4559:data <=32'hFFB50005;
14'd4560:data <=32'hFFC30005;14'd4561:data <=32'hFFCEFFFE;14'd4562:data <=32'hFFD4FFF1;
14'd4563:data <=32'hFFD3FFE5;14'd4564:data <=32'hFFC9FFDA;14'd4565:data <=32'hFFB7FFD4;
14'd4566:data <=32'hFFA4FFD9;14'd4567:data <=32'hFF91FFE7;14'd4568:data <=32'hFF84FFFC;
14'd4569:data <=32'hFF800016;14'd4570:data <=32'hFF860031;14'd4571:data <=32'hFF950047;
14'd4572:data <=32'hFFA90056;14'd4573:data <=32'hFFBF005F;14'd4574:data <=32'hFFD50060;
14'd4575:data <=32'hFFE7005B;14'd4576:data <=32'hFFF70053;14'd4577:data <=32'h00020048;
14'd4578:data <=32'h000A003C;14'd4579:data <=32'h000D002F;14'd4580:data <=32'h000D0021;
14'd4581:data <=32'h00070013;14'd4582:data <=32'hFFFD0009;14'd4583:data <=32'hFFEF0004;
14'd4584:data <=32'hFFDE0005;14'd4585:data <=32'hFFCE000E;14'd4586:data <=32'hFFC2001C;
14'd4587:data <=32'hFFBC0030;14'd4588:data <=32'hFFBD0043;14'd4589:data <=32'hFFC40056;
14'd4590:data <=32'hFFD00065;14'd4591:data <=32'hFFDD0070;14'd4592:data <=32'hFFEA0076;
14'd4593:data <=32'hFFF6007E;14'd4594:data <=32'h00010083;14'd4595:data <=32'h000E008C;
14'd4596:data <=32'h001D0095;14'd4597:data <=32'h0033009F;14'd4598:data <=32'h004D00A4;
14'd4599:data <=32'h006C00A2;14'd4600:data <=32'h008E009C;14'd4601:data <=32'h00AE008A;
14'd4602:data <=32'h00CB0071;14'd4603:data <=32'h00E40052;14'd4604:data <=32'h00F8002D;
14'd4605:data <=32'h01050005;14'd4606:data <=32'h010BFFD9;14'd4607:data <=32'h0109FFAA;
14'd4608:data <=32'h0037FFEE;14'd4609:data <=32'h0053FFEF;14'd4610:data <=32'h007EFFE1;
14'd4611:data <=32'h00E3FF68;14'd4612:data <=32'h00C1FF05;14'd4613:data <=32'h0083FEEC;
14'd4614:data <=32'h0044FEE6;14'd4615:data <=32'h0007FEF0;14'd4616:data <=32'hFFD5FF09;
14'd4617:data <=32'hFFB1FF2B;14'd4618:data <=32'hFF98FF4F;14'd4619:data <=32'hFF8BFF73;
14'd4620:data <=32'hFF85FF95;14'd4621:data <=32'hFF88FFB4;14'd4622:data <=32'hFF90FFCF;
14'd4623:data <=32'hFF9EFFE5;14'd4624:data <=32'hFFAFFFF3;14'd4625:data <=32'hFFC3FFFB;
14'd4626:data <=32'hFFD6FFF9;14'd4627:data <=32'hFFE4FFF1;14'd4628:data <=32'hFFEBFFE3;
14'd4629:data <=32'hFFE9FFD5;14'd4630:data <=32'hFFE0FFCA;14'd4631:data <=32'hFFD2FFC6;
14'd4632:data <=32'hFFC3FFC8;14'd4633:data <=32'hFFB7FFD1;14'd4634:data <=32'hFFB0FFDD;
14'd4635:data <=32'hFFAEFFE9;14'd4636:data <=32'hFFB0FFF4;14'd4637:data <=32'hFFB4FFFB;
14'd4638:data <=32'hFFB60000;14'd4639:data <=32'hFFB70003;14'd4640:data <=32'hFFB70006;
14'd4641:data <=32'hFFB7000B;14'd4642:data <=32'hFFB70012;14'd4643:data <=32'hFFB90018;
14'd4644:data <=32'hFFBD001F;14'd4645:data <=32'hFFC20024;14'd4646:data <=32'hFFC70027;
14'd4647:data <=32'hFFCB0029;14'd4648:data <=32'hFFCF002A;14'd4649:data <=32'hFFD1002C;
14'd4650:data <=32'hFFD4002E;14'd4651:data <=32'hFFD70030;14'd4652:data <=32'hFFDC0031;
14'd4653:data <=32'hFFE0002F;14'd4654:data <=32'hFFE5002B;14'd4655:data <=32'hFFE40024;
14'd4656:data <=32'hFFDE001E;14'd4657:data <=32'hFFD2001A;14'd4658:data <=32'hFFC1001C;
14'd4659:data <=32'hFFAF0029;14'd4660:data <=32'hFF9F003F;14'd4661:data <=32'hFF97005D;
14'd4662:data <=32'hFF9A0083;14'd4663:data <=32'hFFAA00A7;14'd4664:data <=32'hFFC500C9;
14'd4665:data <=32'hFFEB00E4;14'd4666:data <=32'h001800F4;14'd4667:data <=32'h004900FA;
14'd4668:data <=32'h007D00F4;14'd4669:data <=32'h00B000E3;14'd4670:data <=32'h00E100C6;
14'd4671:data <=32'h010C009D;14'd4672:data <=32'h008B0057;14'd4673:data <=32'h00B1004F;
14'd4674:data <=32'h00D1004D;14'd4675:data <=32'h010E005E;14'd4676:data <=32'h011EFFEB;
14'd4677:data <=32'h010AFFB9;14'd4678:data <=32'h00EBFF90;14'd4679:data <=32'h00C7FF72;
14'd4680:data <=32'h00A3FF61;14'd4681:data <=32'h0082FF58;14'd4682:data <=32'h0065FF54;
14'd4683:data <=32'h004AFF53;14'd4684:data <=32'h0032FF54;14'd4685:data <=32'h001AFF58;
14'd4686:data <=32'h0004FF5F;14'd4687:data <=32'hFFF0FF69;14'd4688:data <=32'hFFE0FF76;
14'd4689:data <=32'hFFD4FF86;14'd4690:data <=32'hFFCCFF94;14'd4691:data <=32'hFFC7FFA0;
14'd4692:data <=32'hFFC3FFAA;14'd4693:data <=32'hFFBFFFB4;14'd4694:data <=32'hFFBAFFBE;
14'd4695:data <=32'hFFB6FFCA;14'd4696:data <=32'hFFB4FFD8;14'd4697:data <=32'hFFB6FFE9;
14'd4698:data <=32'hFFBFFFF8;14'd4699:data <=32'hFFCE0002;14'd4700:data <=32'hFFE00006;
14'd4701:data <=32'hFFF00002;14'd4702:data <=32'hFFFEFFF5;14'd4703:data <=32'h0003FFE5;
14'd4704:data <=32'h0001FFD4;14'd4705:data <=32'hFFF8FFC5;14'd4706:data <=32'hFFEAFFBC;
14'd4707:data <=32'hFFD9FFB8;14'd4708:data <=32'hFFC8FFB9;14'd4709:data <=32'hFFB7FFBF;
14'd4710:data <=32'hFFA9FFC9;14'd4711:data <=32'hFF9EFFD5;14'd4712:data <=32'hFF96FFE4;
14'd4713:data <=32'hFF92FFF5;14'd4714:data <=32'hFF910007;14'd4715:data <=32'hFF960018;
14'd4716:data <=32'hFF9F0028;14'd4717:data <=32'hFFAD0032;14'd4718:data <=32'hFFBD0036;
14'd4719:data <=32'hFFCC0032;14'd4720:data <=32'hFFD50029;14'd4721:data <=32'hFFD7001C;
14'd4722:data <=32'hFFD00011;14'd4723:data <=32'hFFC1000A;14'd4724:data <=32'hFFAD000D;
14'd4725:data <=32'hFF9A0019;14'd4726:data <=32'hFF8B002D;14'd4727:data <=32'hFF820049;
14'd4728:data <=32'hFF84006A;14'd4729:data <=32'hFF8E0088;14'd4730:data <=32'hFFA100A5;
14'd4731:data <=32'hFFBA00BC;14'd4732:data <=32'hFFD800CF;14'd4733:data <=32'hFFFA00DD;
14'd4734:data <=32'h002000E4;14'd4735:data <=32'h004A00E3;14'd4736:data <=32'h000D00FC;
14'd4737:data <=32'h004C0113;14'd4738:data <=32'h007C010D;14'd4739:data <=32'h005E00C1;
14'd4740:data <=32'h00810074;14'd4741:data <=32'h00870060;14'd4742:data <=32'h00890051;
14'd4743:data <=32'h00890044;14'd4744:data <=32'h008C003C;14'd4745:data <=32'h00930035;
14'd4746:data <=32'h009F002B;14'd4747:data <=32'h00AE001B;14'd4748:data <=32'h00B90004;
14'd4749:data <=32'h00C0FFE7;14'd4750:data <=32'h00BEFFC7;14'd4751:data <=32'h00B4FFA6;
14'd4752:data <=32'h00A2FF89;14'd4753:data <=32'h008BFF71;14'd4754:data <=32'h0070FF5D;
14'd4755:data <=32'h0052FF51;14'd4756:data <=32'h0031FF48;14'd4757:data <=32'h000EFF47;
14'd4758:data <=32'hFFEAFF4E;14'd4759:data <=32'hFFCAFF5F;14'd4760:data <=32'hFFADFF78;
14'd4761:data <=32'hFF99FF9B;14'd4762:data <=32'hFF93FFC0;14'd4763:data <=32'hFF98FFE5;
14'd4764:data <=32'hFFAA0004;14'd4765:data <=32'hFFC30017;14'd4766:data <=32'hFFE10020;
14'd4767:data <=32'hFFFC001E;14'd4768:data <=32'h00130012;14'd4769:data <=32'h00240000;
14'd4770:data <=32'h002BFFEC;14'd4771:data <=32'h002CFFD8;14'd4772:data <=32'h0029FFC5;
14'd4773:data <=32'h0020FFB5;14'd4774:data <=32'h0014FFA6;14'd4775:data <=32'h0004FF9B;
14'd4776:data <=32'hFFF2FF94;14'd4777:data <=32'hFFDEFF90;14'd4778:data <=32'hFFC9FF92;
14'd4779:data <=32'hFFB6FF99;14'd4780:data <=32'hFFA5FFA5;14'd4781:data <=32'hFF99FFB3;
14'd4782:data <=32'hFF91FFC1;14'd4783:data <=32'hFF8DFFCE;14'd4784:data <=32'hFF89FFD8;
14'd4785:data <=32'hFF85FFE0;14'd4786:data <=32'hFF7FFFE7;14'd4787:data <=32'hFF75FFF1;
14'd4788:data <=32'hFF6B0000;14'd4789:data <=32'hFF610014;14'd4790:data <=32'hFF5C002E;
14'd4791:data <=32'hFF5F004B;14'd4792:data <=32'hFF690068;14'd4793:data <=32'hFF7C0081;
14'd4794:data <=32'hFF930093;14'd4795:data <=32'hFFAD009E;14'd4796:data <=32'hFFC600A5;
14'd4797:data <=32'hFFDD00A6;14'd4798:data <=32'hFFF400A3;14'd4799:data <=32'h0007009E;
14'd4800:data <=32'hFF4C00AE;14'd4801:data <=32'hFF6A00EE;14'd4802:data <=32'hFFA60110;
14'd4803:data <=32'h00170093;14'd4804:data <=32'h002C004C;14'd4805:data <=32'h00210042;
14'd4806:data <=32'h00120040;14'd4807:data <=32'h00060048;14'd4808:data <=32'hFFFF0058;
14'd4809:data <=32'h0003006E;14'd4810:data <=32'h00140083;14'd4811:data <=32'h002D0093;
14'd4812:data <=32'h004F0098;14'd4813:data <=32'h00730091;14'd4814:data <=32'h00950080;
14'd4815:data <=32'h00B00065;14'd4816:data <=32'h00C40044;14'd4817:data <=32'h00CF001F;
14'd4818:data <=32'h00D2FFF9;14'd4819:data <=32'h00CDFFD4;14'd4820:data <=32'h00C0FFAF;
14'd4821:data <=32'h00A9FF8D;14'd4822:data <=32'h008BFF72;14'd4823:data <=32'h0066FF5E;
14'd4824:data <=32'h003DFF57;14'd4825:data <=32'h0014FF5D;14'd4826:data <=32'hFFF1FF6E;
14'd4827:data <=32'hFFD7FF87;14'd4828:data <=32'hFFC9FFA5;14'd4829:data <=32'hFFC5FFC1;
14'd4830:data <=32'hFFCAFFDA;14'd4831:data <=32'hFFD4FFED;14'd4832:data <=32'hFFE0FFF9;
14'd4833:data <=32'hFFED0001;14'd4834:data <=32'hFFFA0005;14'd4835:data <=32'h00060008;
14'd4836:data <=32'h00130007;14'd4837:data <=32'h00200006;14'd4838:data <=32'h002FFFFE;
14'd4839:data <=32'h003BFFF4;14'd4840:data <=32'h0047FFE3;14'd4841:data <=32'h004EFFCF;
14'd4842:data <=32'h004EFFB9;14'd4843:data <=32'h0049FFA2;14'd4844:data <=32'h003EFF8C;
14'd4845:data <=32'h0030FF78;14'd4846:data <=32'h001CFF66;14'd4847:data <=32'h0004FF59;
14'd4848:data <=32'hFFE9FF4C;14'd4849:data <=32'hFFC9FF44;14'd4850:data <=32'hFFA4FF43;
14'd4851:data <=32'hFF7BFF49;14'd4852:data <=32'hFF51FF5B;14'd4853:data <=32'hFF2AFF79;
14'd4854:data <=32'hFF0BFFA4;14'd4855:data <=32'hFEF9FFD7;14'd4856:data <=32'hFEF6000E;
14'd4857:data <=32'hFF000043;14'd4858:data <=32'hFF1A0071;14'd4859:data <=32'hFF3C0095;
14'd4860:data <=32'hFF6300AC;14'd4861:data <=32'hFF8C00B9;14'd4862:data <=32'hFFB200BC;
14'd4863:data <=32'hFFD600B7;14'd4864:data <=32'hFF58002A;14'd4865:data <=32'hFF4E0057;
14'd4866:data <=32'hFF5F0092;14'd4867:data <=32'hFFE000BE;14'd4868:data <=32'h00080074;
14'd4869:data <=32'h000A0060;14'd4870:data <=32'h00050052;14'd4871:data <=32'hFFFB0049;
14'd4872:data <=32'hFFEF004C;14'd4873:data <=32'hFFE70057;14'd4874:data <=32'hFFE80068;
14'd4875:data <=32'hFFF10079;14'd4876:data <=32'h00040086;14'd4877:data <=32'h0019008D;
14'd4878:data <=32'h0032008B;14'd4879:data <=32'h00480084;14'd4880:data <=32'h005C0077;
14'd4881:data <=32'h006B0068;14'd4882:data <=32'h00780058;14'd4883:data <=32'h00820045;
14'd4884:data <=32'h00890031;14'd4885:data <=32'h008E001B;14'd4886:data <=32'h008B0004;
14'd4887:data <=32'h0085FFEE;14'd4888:data <=32'h0079FFDC;14'd4889:data <=32'h0068FFCE;
14'd4890:data <=32'h0057FFC7;14'd4891:data <=32'h0047FFC4;14'd4892:data <=32'h003BFFC6;
14'd4893:data <=32'h0033FFCA;14'd4894:data <=32'h002EFFCB;14'd4895:data <=32'h0028FFCB;
14'd4896:data <=32'h0023FFC9;14'd4897:data <=32'h0019FFC7;14'd4898:data <=32'h000EFFC9;
14'd4899:data <=32'h0002FFD0;14'd4900:data <=32'hFFF9FFDC;14'd4901:data <=32'hFFF5FFEB;
14'd4902:data <=32'hFFF7FFFD;14'd4903:data <=32'h0002000E;14'd4904:data <=32'h00120019;
14'd4905:data <=32'h0028001E;14'd4906:data <=32'h0040001C;14'd4907:data <=32'h00560012;
14'd4908:data <=32'h006A0001;14'd4909:data <=32'h007CFFEB;14'd4910:data <=32'h0087FFCD;
14'd4911:data <=32'h008CFFAB;14'd4912:data <=32'h0089FF86;14'd4913:data <=32'h007BFF5F;
14'd4914:data <=32'h0063FF38;14'd4915:data <=32'h003CFF16;14'd4916:data <=32'h000CFF00;
14'd4917:data <=32'hFFD4FEF7;14'd4918:data <=32'hFF99FEFE;14'd4919:data <=32'hFF64FF16;
14'd4920:data <=32'hFF36FF3B;14'd4921:data <=32'hFF17FF6A;14'd4922:data <=32'hFF05FF9C;
14'd4923:data <=32'hFF01FFCC;14'd4924:data <=32'hFF08FFF9;14'd4925:data <=32'hFF14001F;
14'd4926:data <=32'hFF270040;14'd4927:data <=32'hFF3D005B;14'd4928:data <=32'hFF600027;
14'd4929:data <=32'hFF5B003F;14'd4930:data <=32'hFF52005B;14'd4931:data <=32'hFF2F0078;
14'd4932:data <=32'hFF5B0054;14'd4933:data <=32'hFF680062;14'd4934:data <=32'hFF74006F;
14'd4935:data <=32'hFF80007B;14'd4936:data <=32'hFF8C008B;14'd4937:data <=32'hFF9C009B;
14'd4938:data <=32'hFFB100AC;14'd4939:data <=32'hFFCE00B8;14'd4940:data <=32'hFFEE00BE;
14'd4941:data <=32'h001200BA;14'd4942:data <=32'h003100AB;14'd4943:data <=32'h004B0095;
14'd4944:data <=32'h005A007A;14'd4945:data <=32'h0062005E;14'd4946:data <=32'h00610046;
14'd4947:data <=32'h005B0033;14'd4948:data <=32'h00530023;14'd4949:data <=32'h00490018;
14'd4950:data <=32'h003F0011;14'd4951:data <=32'h0036000D;14'd4952:data <=32'h002B000C;
14'd4953:data <=32'h0021000F;14'd4954:data <=32'h001B0017;14'd4955:data <=32'h001A0020;
14'd4956:data <=32'h001F002B;14'd4957:data <=32'h002A0032;14'd4958:data <=32'h00380034;
14'd4959:data <=32'h0047002E;14'd4960:data <=32'h00540021;14'd4961:data <=32'h005A000F;
14'd4962:data <=32'h0058FFFD;14'd4963:data <=32'h0050FFED;14'd4964:data <=32'h0043FFE3;
14'd4965:data <=32'h0033FFE0;14'd4966:data <=32'h0026FFE4;14'd4967:data <=32'h001CFFED;
14'd4968:data <=32'h0019FFF8;14'd4969:data <=32'h001B0004;14'd4970:data <=32'h0022000E;
14'd4971:data <=32'h002D0015;14'd4972:data <=32'h003B0017;14'd4973:data <=32'h004A0016;
14'd4974:data <=32'h005C0011;14'd4975:data <=32'h006D0007;14'd4976:data <=32'h007DFFF4;
14'd4977:data <=32'h008BFFDD;14'd4978:data <=32'h0091FFBF;14'd4979:data <=32'h0090FF9E;
14'd4980:data <=32'h0084FF7C;14'd4981:data <=32'h006EFF5F;14'd4982:data <=32'h0051FF47;
14'd4983:data <=32'h002EFF3A;14'd4984:data <=32'h000CFF37;14'd4985:data <=32'hFFEEFF39;
14'd4986:data <=32'hFFD4FF42;14'd4987:data <=32'hFFBFFF4B;14'd4988:data <=32'hFFACFF53;
14'd4989:data <=32'hFF9AFF5C;14'd4990:data <=32'hFF87FF65;14'd4991:data <=32'hFF71FF70;
14'd4992:data <=32'hFF2DFFB9;14'd4993:data <=32'hFF1FFFDA;14'd4994:data <=32'hFF22FFEA;
14'd4995:data <=32'hFF3BFF82;14'd4996:data <=32'hFF3AFF67;14'd4997:data <=32'hFF1DFF85;
14'd4998:data <=32'hFF03FFA9;14'd4999:data <=32'hFEF2FFD5;14'd5000:data <=32'hFEE80006;
14'd5001:data <=32'hFEE8003B;14'd5002:data <=32'hFEF70073;14'd5003:data <=32'hFF1500A6;
14'd5004:data <=32'hFF4200D0;14'd5005:data <=32'hFF7800EC;14'd5006:data <=32'hFFB200F6;
14'd5007:data <=32'hFFEA00EF;14'd5008:data <=32'h001900DA;14'd5009:data <=32'h003F00BB;
14'd5010:data <=32'h00570098;14'd5011:data <=32'h00630074;14'd5012:data <=32'h00660052;
14'd5013:data <=32'h00620033;14'd5014:data <=32'h0057001A;14'd5015:data <=32'h00470006;
14'd5016:data <=32'h0033FFF7;14'd5017:data <=32'h001CFFF1;14'd5018:data <=32'h0007FFF3;
14'd5019:data <=32'hFFF3FFFC;14'd5020:data <=32'hFFE6000D;14'd5021:data <=32'hFFE10021;
14'd5022:data <=32'hFFE50035;14'd5023:data <=32'hFFF00043;14'd5024:data <=32'hFFFF004C;
14'd5025:data <=32'h000F004F;14'd5026:data <=32'h001C004C;14'd5027:data <=32'h00250046;
14'd5028:data <=32'h002A0041;14'd5029:data <=32'h002D003E;14'd5030:data <=32'h0030003D;
14'd5031:data <=32'h0036003D;14'd5032:data <=32'h003E003D;14'd5033:data <=32'h0049003C;
14'd5034:data <=32'h00530036;14'd5035:data <=32'h005E002F;14'd5036:data <=32'h00660023;
14'd5037:data <=32'h006C0017;14'd5038:data <=32'h006F000B;14'd5039:data <=32'h0070FFFE;
14'd5040:data <=32'h0072FFF3;14'd5041:data <=32'h0071FFE7;14'd5042:data <=32'h006FFFDA;
14'd5043:data <=32'h006BFFCD;14'd5044:data <=32'h0064FFC1;14'd5045:data <=32'h0059FFB6;
14'd5046:data <=32'h004EFFB0;14'd5047:data <=32'h0042FFAF;14'd5048:data <=32'h003AFFB2;
14'd5049:data <=32'h0039FFB7;14'd5050:data <=32'h003DFFB9;14'd5051:data <=32'h0046FFB6;
14'd5052:data <=32'h0050FFAA;14'd5053:data <=32'h0057FF95;14'd5054:data <=32'h0057FF79;
14'd5055:data <=32'h004BFF5B;14'd5056:data <=32'hFFC5FF33;14'd5057:data <=32'hFFA3FF35;
14'd5058:data <=32'hFF9AFF49;14'd5059:data <=32'h0009FF49;14'd5060:data <=32'h0000FF06;
14'd5061:data <=32'hFFD1FEFE;14'd5062:data <=32'hFF9EFF01;14'd5063:data <=32'hFF6CFF10;
14'd5064:data <=32'hFF3BFF2B;14'd5065:data <=32'hFF11FF54;14'd5066:data <=32'hFEF0FF88;
14'd5067:data <=32'hFEE0FFC5;14'd5068:data <=32'hFEE20002;14'd5069:data <=32'hFEF4003C;
14'd5070:data <=32'hFF13006A;14'd5071:data <=32'hFF3B008C;14'd5072:data <=32'hFF6700A1;
14'd5073:data <=32'hFF9000A9;14'd5074:data <=32'hFFB500A8;14'd5075:data <=32'hFFD400A0;
14'd5076:data <=32'hFFF00094;14'd5077:data <=32'h00070086;14'd5078:data <=32'h00190075;
14'd5079:data <=32'h00270061;14'd5080:data <=32'h002E004C;14'd5081:data <=32'h00300036;
14'd5082:data <=32'h002B0022;14'd5083:data <=32'h00210013;14'd5084:data <=32'h0015000A;
14'd5085:data <=32'h00070006;14'd5086:data <=32'hFFFD0007;14'd5087:data <=32'hFFF50008;
14'd5088:data <=32'hFFED000B;14'd5089:data <=32'hFFE7000F;14'd5090:data <=32'hFFDF0011;
14'd5091:data <=32'hFFD60018;14'd5092:data <=32'hFFCC0023;14'd5093:data <=32'hFFC50033;
14'd5094:data <=32'hFFC10048;14'd5095:data <=32'hFFC70060;14'd5096:data <=32'hFFD40078;
14'd5097:data <=32'hFFEA008D;14'd5098:data <=32'h0007009A;14'd5099:data <=32'h0028009E;
14'd5100:data <=32'h00490099;14'd5101:data <=32'h0067008B;14'd5102:data <=32'h007F0077;
14'd5103:data <=32'h0092005E;14'd5104:data <=32'h009E0043;14'd5105:data <=32'h00A40026;
14'd5106:data <=32'h00A3000B;14'd5107:data <=32'h009EFFF0;14'd5108:data <=32'h0091FFD8;
14'd5109:data <=32'h007EFFC6;14'd5110:data <=32'h0067FFB9;14'd5111:data <=32'h0050FFB8;
14'd5112:data <=32'h003CFFC0;14'd5113:data <=32'h0031FFCE;14'd5114:data <=32'h002FFFDE;
14'd5115:data <=32'h0038FFED;14'd5116:data <=32'h004AFFF4;14'd5117:data <=32'h005FFFF1;
14'd5118:data <=32'h0075FFE2;14'd5119:data <=32'h0084FFC9;14'd5120:data <=32'h0076FFA8;
14'd5121:data <=32'h007AFF88;14'd5122:data <=32'h0069FF7A;14'd5123:data <=32'h004BFFA0;
14'd5124:data <=32'h005DFF5A;14'd5125:data <=32'h0045FF48;14'd5126:data <=32'h0028FF3A;
14'd5127:data <=32'h0009FF32;14'd5128:data <=32'hFFE7FF30;14'd5129:data <=32'hFFC4FF37;
14'd5130:data <=32'hFFA1FF45;14'd5131:data <=32'hFF85FF5D;14'd5132:data <=32'hFF70FF7A;
14'd5133:data <=32'hFF66FF9A;14'd5134:data <=32'hFF64FFB7;14'd5135:data <=32'hFF68FFCF;
14'd5136:data <=32'hFF6FFFE0;14'd5137:data <=32'hFF75FFEE;14'd5138:data <=32'hFF79FFF9;
14'd5139:data <=32'hFF790004;14'd5140:data <=32'hFF7A0013;14'd5141:data <=32'hFF7E0024;
14'd5142:data <=32'hFF860036;14'd5143:data <=32'hFF930046;14'd5144:data <=32'hFFA30052;
14'd5145:data <=32'hFFB7005A;14'd5146:data <=32'hFFCB005C;14'd5147:data <=32'hFFDD005B;
14'd5148:data <=32'hFFED0056;14'd5149:data <=32'hFFFC004F;14'd5150:data <=32'h00090045;
14'd5151:data <=32'h00130037;14'd5152:data <=32'h001B0026;14'd5153:data <=32'h001C0011;
14'd5154:data <=32'h0015FFFC;14'd5155:data <=32'h0006FFE9;14'd5156:data <=32'hFFEFFFDC;
14'd5157:data <=32'hFFD3FFDA;14'd5158:data <=32'hFFB6FFE3;14'd5159:data <=32'hFF9CFFF6;
14'd5160:data <=32'hFF8B0013;14'd5161:data <=32'hFF840036;14'd5162:data <=32'hFF880059;
14'd5163:data <=32'hFF98007A;14'd5164:data <=32'hFFAF0093;14'd5165:data <=32'hFFCB00A6;
14'd5166:data <=32'hFFEA00B1;14'd5167:data <=32'h000900B5;14'd5168:data <=32'h002800B3;
14'd5169:data <=32'h004500AA;14'd5170:data <=32'h005F009D;14'd5171:data <=32'h00760089;
14'd5172:data <=32'h00870072;14'd5173:data <=32'h00920059;14'd5174:data <=32'h00950040;
14'd5175:data <=32'h0092002B;14'd5176:data <=32'h008C001B;14'd5177:data <=32'h00850010;
14'd5178:data <=32'h0082000C;14'd5179:data <=32'h00840009;14'd5180:data <=32'h008A0004;
14'd5181:data <=32'h0093FFF9;14'd5182:data <=32'h009DFFE8;14'd5183:data <=32'h00A2FFD1;
14'd5184:data <=32'h00470035;14'd5185:data <=32'h006F0031;14'd5186:data <=32'h00890013;
14'd5187:data <=32'h0072FF96;14'd5188:data <=32'h0079FF57;14'd5189:data <=32'h0057FF4E;
14'd5190:data <=32'h0037FF4D;14'd5191:data <=32'h001AFF53;14'd5192:data <=32'h0001FF5B;
14'd5193:data <=32'hFFEAFF69;14'd5194:data <=32'hFFD8FF7A;14'd5195:data <=32'hFFCCFF8E;
14'd5196:data <=32'hFFC8FFA4;14'd5197:data <=32'hFFCBFFB8;14'd5198:data <=32'hFFD5FFC6;
14'd5199:data <=32'hFFE3FFCA;14'd5200:data <=32'hFFEFFFC7;14'd5201:data <=32'hFFF6FFBA;
14'd5202:data <=32'hFFF3FFAB;14'd5203:data <=32'hFFE6FF9D;14'd5204:data <=32'hFFD3FF95;
14'd5205:data <=32'hFFBCFF95;14'd5206:data <=32'hFFA5FF9E;14'd5207:data <=32'hFF91FFAE;
14'd5208:data <=32'hFF84FFC3;14'd5209:data <=32'hFF7DFFDA;14'd5210:data <=32'hFF7BFFF2;
14'd5211:data <=32'hFF7F0008;14'd5212:data <=32'hFF87001D;14'd5213:data <=32'hFF950030;
14'd5214:data <=32'hFFA7003F;14'd5215:data <=32'hFFBC0049;14'd5216:data <=32'hFFD4004A;
14'd5217:data <=32'hFFEC0044;14'd5218:data <=32'h00000036;14'd5219:data <=32'h000B0022;
14'd5220:data <=32'h000D000B;14'd5221:data <=32'h0006FFF4;14'd5222:data <=32'hFFF6FFE4;
14'd5223:data <=32'hFFE2FFDC;14'd5224:data <=32'hFFCCFFDC;14'd5225:data <=32'hFFB9FFE4;
14'd5226:data <=32'hFFA9FFF0;14'd5227:data <=32'hFF9F0000;14'd5228:data <=32'hFF980010;
14'd5229:data <=32'hFF950021;14'd5230:data <=32'hFF930031;14'd5231:data <=32'hFF930040;
14'd5232:data <=32'hFF940053;14'd5233:data <=32'hFF980067;14'd5234:data <=32'hFFA1007C;
14'd5235:data <=32'hFFAE0091;14'd5236:data <=32'hFFC100A4;14'd5237:data <=32'hFFD600B2;
14'd5238:data <=32'hFFEF00BE;14'd5239:data <=32'h000900C5;14'd5240:data <=32'h002400CA;
14'd5241:data <=32'h004200CD;14'd5242:data <=32'h006200CB;14'd5243:data <=32'h008600C5;
14'd5244:data <=32'h00AD00B6;14'd5245:data <=32'h00D4009D;14'd5246:data <=32'h00F50077;
14'd5247:data <=32'h010E0047;14'd5248:data <=32'h00260031;14'd5249:data <=32'h00400044;
14'd5250:data <=32'h006E004B;14'd5251:data <=32'h00F9FFF8;14'd5252:data <=32'h0106FF99;
14'd5253:data <=32'h00E1FF71;14'd5254:data <=32'h00B6FF55;14'd5255:data <=32'h0089FF46;
14'd5256:data <=32'h005FFF41;14'd5257:data <=32'h0035FF45;14'd5258:data <=32'h0010FF53;
14'd5259:data <=32'hFFF1FF68;14'd5260:data <=32'hFFDDFF84;14'd5261:data <=32'hFFD4FFA3;
14'd5262:data <=32'hFFD8FFBF;14'd5263:data <=32'hFFE5FFD4;14'd5264:data <=32'hFFF7FFE0;
14'd5265:data <=32'h0009FFDE;14'd5266:data <=32'h0017FFD4;14'd5267:data <=32'h001DFFC6;
14'd5268:data <=32'h001AFFB6;14'd5269:data <=32'h0012FFA8;14'd5270:data <=32'h0004FFA0;
14'd5271:data <=32'hFFF4FF9D;14'd5272:data <=32'hFFE6FF9E;14'd5273:data <=32'hFFD9FFA3;
14'd5274:data <=32'hFFCDFFA8;14'd5275:data <=32'hFFC4FFAF;14'd5276:data <=32'hFFB9FFB9;
14'd5277:data <=32'hFFB2FFC3;14'd5278:data <=32'hFFADFFD1;14'd5279:data <=32'hFFABFFE0;
14'd5280:data <=32'hFFAEFFEC;14'd5281:data <=32'hFFB5FFF7;14'd5282:data <=32'hFFBDFFFF;
14'd5283:data <=32'hFFC60001;14'd5284:data <=32'hFFCD0000;14'd5285:data <=32'hFFD1FFFD;
14'd5286:data <=32'hFFD1FFFB;14'd5287:data <=32'hFFCEFFFA;14'd5288:data <=32'hFFCDFFFC;
14'd5289:data <=32'hFFCC0000;14'd5290:data <=32'hFFCF0003;14'd5291:data <=32'hFFD40003;
14'd5292:data <=32'hFFD90000;14'd5293:data <=32'hFFDCFFF7;14'd5294:data <=32'hFFD8FFED;
14'd5295:data <=32'hFFCFFFE3;14'd5296:data <=32'hFFBEFFDA;14'd5297:data <=32'hFFA9FFD9;
14'd5298:data <=32'hFF8FFFDF;14'd5299:data <=32'hFF78FFEE;14'd5300:data <=32'hFF630006;
14'd5301:data <=32'hFF540024;14'd5302:data <=32'hFF4B0046;14'd5303:data <=32'hFF4A006E;
14'd5304:data <=32'hFF510097;14'd5305:data <=32'hFF6200C2;14'd5306:data <=32'hFF7F00EB;
14'd5307:data <=32'hFFA80111;14'd5308:data <=32'hFFDE012E;14'd5309:data <=32'h001E013B;
14'd5310:data <=32'h00620137;14'd5311:data <=32'h00A4011F;14'd5312:data <=32'h003B008D;
14'd5313:data <=32'h00590099;14'd5314:data <=32'h007200AD;14'd5315:data <=32'h00B400DD;
14'd5316:data <=32'h00F10081;14'd5317:data <=32'h00F70052;14'd5318:data <=32'h00F40027;
14'd5319:data <=32'h00EA0002;14'd5320:data <=32'h00DBFFDF;14'd5321:data <=32'h00C7FFC1;
14'd5322:data <=32'h00AEFFAA;14'd5323:data <=32'h0093FF9A;14'd5324:data <=32'h0077FF91;
14'd5325:data <=32'h005EFF91;14'd5326:data <=32'h004AFF96;14'd5327:data <=32'h003EFF9C;
14'd5328:data <=32'h0035FFA1;14'd5329:data <=32'h0030FFA3;14'd5330:data <=32'h002AFFA1;
14'd5331:data <=32'h0021FF9E;14'd5332:data <=32'h0015FF9B;14'd5333:data <=32'h0006FF9C;
14'd5334:data <=32'hFFF7FFA3;14'd5335:data <=32'hFFECFFAF;14'd5336:data <=32'hFFE6FFBE;
14'd5337:data <=32'hFFE6FFCC;14'd5338:data <=32'hFFEBFFD7;14'd5339:data <=32'hFFF3FFDD;
14'd5340:data <=32'hFFFBFFDF;14'd5341:data <=32'h0001FFDC;14'd5342:data <=32'h0007FFD7;
14'd5343:data <=32'h0009FFD3;14'd5344:data <=32'h0009FFCB;14'd5345:data <=32'h0007FFC4;
14'd5346:data <=32'h0004FFBD;14'd5347:data <=32'hFFFEFFB5;14'd5348:data <=32'hFFF5FFAD;
14'd5349:data <=32'hFFE7FFA9;14'd5350:data <=32'hFFD6FFA7;14'd5351:data <=32'hFFC5FFAD;
14'd5352:data <=32'hFFB5FFB9;14'd5353:data <=32'hFFABFFCA;14'd5354:data <=32'hFFA9FFDD;
14'd5355:data <=32'hFFAEFFEE;14'd5356:data <=32'hFFBAFFFB;14'd5357:data <=32'hFFC9FFFF;
14'd5358:data <=32'hFFD8FFFC;14'd5359:data <=32'hFFE1FFF1;14'd5360:data <=32'hFFE3FFE1;
14'd5361:data <=32'hFFDCFFD1;14'd5362:data <=32'hFFCEFFC5;14'd5363:data <=32'hFFBBFFBD;
14'd5364:data <=32'hFFA3FFBB;14'd5365:data <=32'hFF8AFFC1;14'd5366:data <=32'hFF71FFCE;
14'd5367:data <=32'hFF5AFFE2;14'd5368:data <=32'hFF45FFFC;14'd5369:data <=32'hFF35001E;
14'd5370:data <=32'hFF2D0047;14'd5371:data <=32'hFF310075;14'd5372:data <=32'hFF4100A3;
14'd5373:data <=32'hFF5E00CE;14'd5374:data <=32'hFF8800EF;14'd5375:data <=32'hFFB90104;
14'd5376:data <=32'hFF9300E6;14'd5377:data <=32'hFFBC0110;14'd5378:data <=32'hFFDE011F;
14'd5379:data <=32'hFFD300E3;14'd5380:data <=32'h001200B4;14'd5381:data <=32'h002100AF;
14'd5382:data <=32'h003200AC;14'd5383:data <=32'h004400A8;14'd5384:data <=32'h005800A4;
14'd5385:data <=32'h006D009B;14'd5386:data <=32'h0083008C;14'd5387:data <=32'h0096007A;
14'd5388:data <=32'h00A50065;14'd5389:data <=32'h00B2004E;14'd5390:data <=32'h00BB0036;
14'd5391:data <=32'h00C2001B;14'd5392:data <=32'h00C7FFFE;14'd5393:data <=32'h00C6FFDC;
14'd5394:data <=32'h00BDFFBA;14'd5395:data <=32'h00AAFF98;14'd5396:data <=32'h008CFF7B;
14'd5397:data <=32'h0067FF67;14'd5398:data <=32'h003EFF61;14'd5399:data <=32'h0015FF67;
14'd5400:data <=32'hFFF5FF79;14'd5401:data <=32'hFFDCFF93;14'd5402:data <=32'hFFCFFFB0;
14'd5403:data <=32'hFFCDFFCD;14'd5404:data <=32'hFFD2FFE6;14'd5405:data <=32'hFFDFFFFA;
14'd5406:data <=32'hFFEF0007;14'd5407:data <=32'h0000000F;14'd5408:data <=32'h00130011;
14'd5409:data <=32'h0026000C;14'd5410:data <=32'h00370003;14'd5411:data <=32'h0045FFF3;
14'd5412:data <=32'h004CFFDE;14'd5413:data <=32'h004EFFC7;14'd5414:data <=32'h0047FFB0;
14'd5415:data <=32'h0038FF9D;14'd5416:data <=32'h0025FF91;14'd5417:data <=32'h000FFF8C;
14'd5418:data <=32'hFFFDFF8D;14'd5419:data <=32'hFFEEFF93;14'd5420:data <=32'hFFE3FF9A;
14'd5421:data <=32'hFFDEFFA0;14'd5422:data <=32'hFFDBFFA3;14'd5423:data <=32'hFFD6FFA2;
14'd5424:data <=32'hFFCFFF9E;14'd5425:data <=32'hFFC4FF9C;14'd5426:data <=32'hFFB5FF9B;
14'd5427:data <=32'hFFA4FF9F;14'd5428:data <=32'hFF93FFA7;14'd5429:data <=32'hFF84FFB3;
14'd5430:data <=32'hFF76FFC2;14'd5431:data <=32'hFF6DFFD3;14'd5432:data <=32'hFF65FFE6;
14'd5433:data <=32'hFF5EFFF9;14'd5434:data <=32'hFF5B000E;14'd5435:data <=32'hFF5A0026;
14'd5436:data <=32'hFF60003F;14'd5437:data <=32'hFF6B0057;14'd5438:data <=32'hFF7C006B;
14'd5439:data <=32'hFF930078;14'd5440:data <=32'hFEFB0048;14'd5441:data <=32'hFEFC008A;
14'd5442:data <=32'hFF1E00B8;14'd5443:data <=32'hFFA10068;14'd5444:data <=32'hFFC60039;
14'd5445:data <=32'hFFB9003A;14'd5446:data <=32'hFFAC0044;14'd5447:data <=32'hFFA20058;
14'd5448:data <=32'hFFA20071;14'd5449:data <=32'hFFA9008C;14'd5450:data <=32'hFFBC00A5;
14'd5451:data <=32'hFFD400B8;14'd5452:data <=32'hFFF200C8;14'd5453:data <=32'h001500D1;
14'd5454:data <=32'h003B00D2;14'd5455:data <=32'h006200CC;14'd5456:data <=32'h008B00BB;
14'd5457:data <=32'h00B0009F;14'd5458:data <=32'h00CE0077;14'd5459:data <=32'h00E00049;
14'd5460:data <=32'h00E40016;14'd5461:data <=32'h00D8FFE4;14'd5462:data <=32'h00BFFFBA;
14'd5463:data <=32'h009CFF9D;14'd5464:data <=32'h0076FF8B;14'd5465:data <=32'h0051FF87;
14'd5466:data <=32'h002FFF8D;14'd5467:data <=32'h0015FF99;14'd5468:data <=32'h0001FFA9;
14'd5469:data <=32'hFFF3FFBB;14'd5470:data <=32'hFFE9FFCE;14'd5471:data <=32'hFFE5FFE1;
14'd5472:data <=32'hFFE7FFF5;14'd5473:data <=32'hFFEE0007;14'd5474:data <=32'hFFF90016;
14'd5475:data <=32'h00090022;14'd5476:data <=32'h001D0026;14'd5477:data <=32'h00310025;
14'd5478:data <=32'h0044001D;14'd5479:data <=32'h00530012;14'd5480:data <=32'h005E0002;
14'd5481:data <=32'h0065FFF3;14'd5482:data <=32'h006AFFE3;14'd5483:data <=32'h006FFFD2;
14'd5484:data <=32'h0071FFC0;14'd5485:data <=32'h0074FFAA;14'd5486:data <=32'h0071FF90;
14'd5487:data <=32'h0067FF74;14'd5488:data <=32'h0055FF56;14'd5489:data <=32'h0039FF3C;
14'd5490:data <=32'h0014FF29;14'd5491:data <=32'hFFE9FF1F;14'd5492:data <=32'hFFBCFF22;
14'd5493:data <=32'hFF91FF31;14'd5494:data <=32'hFF6DFF4B;14'd5495:data <=32'hFF50FF69;
14'd5496:data <=32'hFF3CFF8D;14'd5497:data <=32'hFF30FFB3;14'd5498:data <=32'hFF2CFFD9;
14'd5499:data <=32'hFF31FFFE;14'd5500:data <=32'hFF3D0020;14'd5501:data <=32'hFF51003F;
14'd5502:data <=32'hFF6C0055;14'd5503:data <=32'hFF8B0062;14'd5504:data <=32'hFF50FFB7;
14'd5505:data <=32'hFF31FFD6;14'd5506:data <=32'hFF28000A;14'd5507:data <=32'hFF92005B;
14'd5508:data <=32'hFFC50025;14'd5509:data <=32'hFFBF0018;14'd5510:data <=32'hFFB20014;
14'd5511:data <=32'hFFA20017;14'd5512:data <=32'hFF960024;14'd5513:data <=32'hFF8E0037;
14'd5514:data <=32'hFF8C004B;14'd5515:data <=32'hFF910061;14'd5516:data <=32'hFF9A0076;
14'd5517:data <=32'hFFA8008A;14'd5518:data <=32'hFFBA009C;14'd5519:data <=32'hFFD300AB;
14'd5520:data <=32'hFFF000B6;14'd5521:data <=32'h001100B9;14'd5522:data <=32'h003400B3;
14'd5523:data <=32'h005300A3;14'd5524:data <=32'h006D008A;14'd5525:data <=32'h007D006D;
14'd5526:data <=32'h0083004F;14'd5527:data <=32'h00810034;14'd5528:data <=32'h0079001E;
14'd5529:data <=32'h0070000E;14'd5530:data <=32'h00650004;14'd5531:data <=32'h005EFFFA;
14'd5532:data <=32'h0057FFF2;14'd5533:data <=32'h004FFFE9;14'd5534:data <=32'h0046FFE1;
14'd5535:data <=32'h003AFFDA;14'd5536:data <=32'h002CFFD7;14'd5537:data <=32'h001CFFD8;
14'd5538:data <=32'h000EFFDF;14'd5539:data <=32'h0003FFEA;14'd5540:data <=32'hFFFCFFF8;
14'd5541:data <=32'hFFFA0007;14'd5542:data <=32'hFFFD0016;14'd5543:data <=32'h00030024;
14'd5544:data <=32'h000D0031;14'd5545:data <=32'h001C003E;14'd5546:data <=32'h00300047;
14'd5547:data <=32'h004A004D;14'd5548:data <=32'h0066004B;14'd5549:data <=32'h00870041;
14'd5550:data <=32'h00A7002A;14'd5551:data <=32'h00C20008;14'd5552:data <=32'h00D3FFDA;
14'd5553:data <=32'h00D6FFA8;14'd5554:data <=32'h00CAFF74;14'd5555:data <=32'h00AEFF45;
14'd5556:data <=32'h0087FF1E;14'd5557:data <=32'h0057FF05;14'd5558:data <=32'h0025FEF9;
14'd5559:data <=32'hFFF3FEF8;14'd5560:data <=32'hFFC3FF03;14'd5561:data <=32'hFF99FF17;
14'd5562:data <=32'hFF75FF31;14'd5563:data <=32'hFF58FF51;14'd5564:data <=32'hFF43FF79;
14'd5565:data <=32'hFF39FFA0;14'd5566:data <=32'hFF39FFC9;14'd5567:data <=32'hFF44FFEC;
14'd5568:data <=32'hFF85FFC5;14'd5569:data <=32'hFF7BFFCE;14'd5570:data <=32'hFF65FFD9;
14'd5571:data <=32'hFF37FFEE;14'd5572:data <=32'hFF66FFD5;14'd5573:data <=32'hFF60FFE1;
14'd5574:data <=32'hFF59FFF1;14'd5575:data <=32'hFF510005;14'd5576:data <=32'hFF510020;
14'd5577:data <=32'hFF57003A;14'd5578:data <=32'hFF640054;14'd5579:data <=32'hFF770068;
14'd5580:data <=32'hFF8E0076;14'd5581:data <=32'hFFA4007F;14'd5582:data <=32'hFFBA0083;
14'd5583:data <=32'hFFCE0084;14'd5584:data <=32'hFFE10082;14'd5585:data <=32'hFFF3007D;
14'd5586:data <=32'h00050075;14'd5587:data <=32'h00130068;14'd5588:data <=32'h001D0059;
14'd5589:data <=32'h00200049;14'd5590:data <=32'h001C003A;14'd5591:data <=32'h00150031;
14'd5592:data <=32'h000B002F;14'd5593:data <=32'h00020034;14'd5594:data <=32'h0000003D;
14'd5595:data <=32'h00050049;14'd5596:data <=32'h00100050;14'd5597:data <=32'h001F0052;
14'd5598:data <=32'h002F004E;14'd5599:data <=32'h003B0045;14'd5600:data <=32'h00430036;
14'd5601:data <=32'h00460027;14'd5602:data <=32'h00430019;14'd5603:data <=32'h003C000D;
14'd5604:data <=32'h00340005;14'd5605:data <=32'h00290001;14'd5606:data <=32'h001E0001;
14'd5607:data <=32'h00130003;14'd5608:data <=32'h000A000B;14'd5609:data <=32'h00020018;
14'd5610:data <=32'hFFFF0028;14'd5611:data <=32'h0004003C;14'd5612:data <=32'h00100050;
14'd5613:data <=32'h00270060;14'd5614:data <=32'h00430068;14'd5615:data <=32'h00660067;
14'd5616:data <=32'h00880059;14'd5617:data <=32'h00A50041;14'd5618:data <=32'h00B90021;
14'd5619:data <=32'h00C4FFFB;14'd5620:data <=32'h00C4FFD5;14'd5621:data <=32'h00BDFFB3;
14'd5622:data <=32'h00AEFF96;14'd5623:data <=32'h009DFF7D;14'd5624:data <=32'h0089FF66;
14'd5625:data <=32'h0073FF55;14'd5626:data <=32'h005AFF44;14'd5627:data <=32'h003FFF38;
14'd5628:data <=32'h0023FF31;14'd5629:data <=32'h0007FF2F;14'd5630:data <=32'hFFEAFF32;
14'd5631:data <=32'hFFD1FF3A;14'd5632:data <=32'hFF82FF7A;14'd5633:data <=32'hFF78FF8D;
14'd5634:data <=32'hFF7CFF8E;14'd5635:data <=32'hFFAAFF2B;14'd5636:data <=32'hFFB3FF08;
14'd5637:data <=32'hFF84FF0F;14'd5638:data <=32'hFF55FF24;14'd5639:data <=32'hFF28FF44;
14'd5640:data <=32'hFF06FF72;14'd5641:data <=32'hFEF1FFAA;14'd5642:data <=32'hFEEDFFE4;
14'd5643:data <=32'hFEF8001B;14'd5644:data <=32'hFF0F004A;14'd5645:data <=32'hFF30006F;
14'd5646:data <=32'hFF56008B;14'd5647:data <=32'hFF7E009A;14'd5648:data <=32'hFFA600A1;
14'd5649:data <=32'hFFCC009E;14'd5650:data <=32'hFFEE0094;14'd5651:data <=32'h000C0080;
14'd5652:data <=32'h00200066;14'd5653:data <=32'h002C0048;14'd5654:data <=32'h002B002A;
14'd5655:data <=32'h001F0011;14'd5656:data <=32'h000CFFFF;14'd5657:data <=32'hFFF5FFFA;
14'd5658:data <=32'hFFE2FFFF;14'd5659:data <=32'hFFD2000B;14'd5660:data <=32'hFFCA001B;
14'd5661:data <=32'hFFCB002C;14'd5662:data <=32'hFFD0003A;14'd5663:data <=32'hFFD90043;
14'd5664:data <=32'hFFE30048;14'd5665:data <=32'hFFEC004B;14'd5666:data <=32'hFFF4004C;
14'd5667:data <=32'hFFFB004C;14'd5668:data <=32'h0001004D;14'd5669:data <=32'h0008004C;
14'd5670:data <=32'h000F004B;14'd5671:data <=32'h0014004A;14'd5672:data <=32'h00180046;
14'd5673:data <=32'h001B0043;14'd5674:data <=32'h001D0043;14'd5675:data <=32'h001F0044;
14'd5676:data <=32'h00220048;14'd5677:data <=32'h0028004C;14'd5678:data <=32'h00330051;
14'd5679:data <=32'h00420051;14'd5680:data <=32'h004F004B;14'd5681:data <=32'h005C0042;
14'd5682:data <=32'h00660034;14'd5683:data <=32'h006A0026;14'd5684:data <=32'h0069001A;
14'd5685:data <=32'h00660012;14'd5686:data <=32'h0063000F;14'd5687:data <=32'h00660010;
14'd5688:data <=32'h006C0010;14'd5689:data <=32'h0077000E;14'd5690:data <=32'h00870006;
14'd5691:data <=32'h0096FFF8;14'd5692:data <=32'h00A4FFE3;14'd5693:data <=32'h00ADFFC9;
14'd5694:data <=32'h00B1FFAC;14'd5695:data <=32'h00AEFF8C;14'd5696:data <=32'h0029FF46;
14'd5697:data <=32'h0018FF41;14'd5698:data <=32'h0017FF4D;14'd5699:data <=32'h008FFF5F;
14'd5700:data <=32'h00A3FF12;14'd5701:data <=32'h0075FEEA;14'd5702:data <=32'h003AFED0;
14'd5703:data <=32'hFFF9FEC4;14'd5704:data <=32'hFFB6FECD;14'd5705:data <=32'hFF79FEE8;
14'd5706:data <=32'hFF49FF12;14'd5707:data <=32'hFF26FF44;14'd5708:data <=32'hFF13FF78;
14'd5709:data <=32'hFF0DFFAC;14'd5710:data <=32'hFF11FFDC;14'd5711:data <=32'hFF1E0007;
14'd5712:data <=32'hFF33002B;14'd5713:data <=32'hFF4E004A;14'd5714:data <=32'hFF6D0061;
14'd5715:data <=32'hFF90006E;14'd5716:data <=32'hFFB20071;14'd5717:data <=32'hFFD2006A;
14'd5718:data <=32'hFFEA005B;14'd5719:data <=32'hFFFA0048;14'd5720:data <=32'h00010034;
14'd5721:data <=32'h00010024;14'd5722:data <=32'hFFFC0017;14'd5723:data <=32'hFFF60010;
14'd5724:data <=32'hFFF1000D;14'd5725:data <=32'hFFEE000A;14'd5726:data <=32'hFFEB0007;
14'd5727:data <=32'hFFE80003;14'd5728:data <=32'hFFE2FFFE;14'd5729:data <=32'hFFD8FFFA;
14'd5730:data <=32'hFFCBFFFB;14'd5731:data <=32'hFFBD0001;14'd5732:data <=32'hFFB0000B;
14'd5733:data <=32'hFFA7001D;14'd5734:data <=32'hFFA30030;14'd5735:data <=32'hFFA50045;
14'd5736:data <=32'hFFAC0059;14'd5737:data <=32'hFFB7006A;14'd5738:data <=32'hFFC7007A;
14'd5739:data <=32'hFFD80086;14'd5740:data <=32'hFFEE008F;14'd5741:data <=32'h00050095;
14'd5742:data <=32'h001D0095;14'd5743:data <=32'h0039008E;14'd5744:data <=32'h00500080;
14'd5745:data <=32'h0064006C;14'd5746:data <=32'h006F0052;14'd5747:data <=32'h00700038;
14'd5748:data <=32'h00680021;14'd5749:data <=32'h00580012;14'd5750:data <=32'h0047000D;
14'd5751:data <=32'h00370010;14'd5752:data <=32'h002C001D;14'd5753:data <=32'h002C002D;
14'd5754:data <=32'h0035003D;14'd5755:data <=32'h00460049;14'd5756:data <=32'h005D004E;
14'd5757:data <=32'h0076004D;14'd5758:data <=32'h00910043;14'd5759:data <=32'h00AB0031;
14'd5760:data <=32'h0098FFFC;14'd5761:data <=32'h00B0FFE8;14'd5762:data <=32'h00B1FFDD;
14'd5763:data <=32'h00A0FFFF;14'd5764:data <=32'h00D6FFB9;14'd5765:data <=32'h00CEFF8F;
14'd5766:data <=32'h00B7FF66;14'd5767:data <=32'h0098FF44;14'd5768:data <=32'h006FFF2D;
14'd5769:data <=32'h0045FF24;14'd5770:data <=32'h001CFF26;14'd5771:data <=32'hFFF9FF2F;
14'd5772:data <=32'hFFDEFF3D;14'd5773:data <=32'hFFC8FF4C;14'd5774:data <=32'hFFB6FF5C;
14'd5775:data <=32'hFFA6FF6C;14'd5776:data <=32'hFF96FF7D;14'd5777:data <=32'hFF8AFF90;
14'd5778:data <=32'hFF81FFA4;14'd5779:data <=32'hFF7DFFBB;14'd5780:data <=32'hFF7CFFD0;
14'd5781:data <=32'hFF81FFE3;14'd5782:data <=32'hFF86FFF3;14'd5783:data <=32'hFF8D0001;
14'd5784:data <=32'hFF94000D;14'd5785:data <=32'hFF9B0019;14'd5786:data <=32'hFFA40025;
14'd5787:data <=32'hFFB10031;14'd5788:data <=32'hFFC2003B;14'd5789:data <=32'hFFD6003E;
14'd5790:data <=32'hFFEC003B;14'd5791:data <=32'h0002002F;14'd5792:data <=32'h0010001C;
14'd5793:data <=32'h00160003;14'd5794:data <=32'h0011FFE9;14'd5795:data <=32'h0003FFD4;
14'd5796:data <=32'hFFECFFC4;14'd5797:data <=32'hFFD3FFBF;14'd5798:data <=32'hFFB8FFC2;
14'd5799:data <=32'hFF9EFFCC;14'd5800:data <=32'hFF89FFDE;14'd5801:data <=32'hFF79FFF6;
14'd5802:data <=32'hFF6F0011;14'd5803:data <=32'hFF6B002E;14'd5804:data <=32'hFF6F004D;
14'd5805:data <=32'hFF79006B;14'd5806:data <=32'hFF8D0087;14'd5807:data <=32'hFFA6009C;
14'd5808:data <=32'hFFC600AB;14'd5809:data <=32'hFFE700AE;14'd5810:data <=32'h000700A8;
14'd5811:data <=32'h0020009B;14'd5812:data <=32'h00310089;14'd5813:data <=32'h00390077;
14'd5814:data <=32'h003A0069;14'd5815:data <=32'h00380061;14'd5816:data <=32'h0037005F;
14'd5817:data <=32'h003A0061;14'd5818:data <=32'h00410065;14'd5819:data <=32'h004E0067;
14'd5820:data <=32'h005C0066;14'd5821:data <=32'h006D0061;14'd5822:data <=32'h007D0057;
14'd5823:data <=32'h008C004B;14'd5824:data <=32'h001B0079;14'd5825:data <=32'h00460092;
14'd5826:data <=32'h0070008B;14'd5827:data <=32'h00890019;14'd5828:data <=32'h00BBFFE2;
14'd5829:data <=32'h00AEFFC6;14'd5830:data <=32'h009BFFAD;14'd5831:data <=32'h0084FF9A;
14'd5832:data <=32'h0069FF91;14'd5833:data <=32'h004EFF90;14'd5834:data <=32'h003AFF99;
14'd5835:data <=32'h002EFFA6;14'd5836:data <=32'h0029FFB1;14'd5837:data <=32'h002DFFB9;
14'd5838:data <=32'h0033FFB9;14'd5839:data <=32'h0039FFB3;14'd5840:data <=32'h003AFFA7;
14'd5841:data <=32'h0036FF99;14'd5842:data <=32'h002CFF8B;14'd5843:data <=32'h001EFF7F;
14'd5844:data <=32'h000CFF78;14'd5845:data <=32'hFFF7FF74;14'd5846:data <=32'hFFE3FF73;
14'd5847:data <=32'hFFCDFF76;14'd5848:data <=32'hFFB4FF7F;14'd5849:data <=32'hFF9EFF8F;
14'd5850:data <=32'hFF8BFFA5;14'd5851:data <=32'hFF7FFFC3;14'd5852:data <=32'hFF7CFFE2;
14'd5853:data <=32'hFF850002;14'd5854:data <=32'hFF97001C;14'd5855:data <=32'hFFB1002E;
14'd5856:data <=32'hFFCE0033;14'd5857:data <=32'hFFE8002E;14'd5858:data <=32'hFFFE001F;
14'd5859:data <=32'h000C000C;14'd5860:data <=32'h0010FFF7;14'd5861:data <=32'h000DFFE3;
14'd5862:data <=32'h0004FFD2;14'd5863:data <=32'hFFF7FFC5;14'd5864:data <=32'hFFE7FFBC;
14'd5865:data <=32'hFFD6FFB6;14'd5866:data <=32'hFFC3FFB5;14'd5867:data <=32'hFFADFFB8;
14'd5868:data <=32'hFF99FFC0;14'd5869:data <=32'hFF86FFCE;14'd5870:data <=32'hFF76FFE0;
14'd5871:data <=32'hFF6AFFF7;14'd5872:data <=32'hFF650010;14'd5873:data <=32'hFF650028;
14'd5874:data <=32'hFF6A003E;14'd5875:data <=32'hFF710052;14'd5876:data <=32'hFF780063;
14'd5877:data <=32'hFF7E0075;14'd5878:data <=32'hFF860088;14'd5879:data <=32'hFF91009E;
14'd5880:data <=32'hFFA100B8;14'd5881:data <=32'hFFBA00D1;14'd5882:data <=32'hFFDC00E6;
14'd5883:data <=32'h000400F1;14'd5884:data <=32'h003100F2;14'd5885:data <=32'h005C00E9;
14'd5886:data <=32'h008600D3;14'd5887:data <=32'h00A700B7;14'd5888:data <=32'hFFD6004C;
14'd5889:data <=32'hFFE10079;14'd5890:data <=32'h000C009F;14'd5891:data <=32'h00B60084;
14'd5892:data <=32'h00F2003B;14'd5893:data <=32'h00EB000A;14'd5894:data <=32'h00D8FFDE;
14'd5895:data <=32'h00BCFFBA;14'd5896:data <=32'h0097FFA2;14'd5897:data <=32'h006FFF99;
14'd5898:data <=32'h004BFF9E;14'd5899:data <=32'h002FFFAE;14'd5900:data <=32'h0020FFC3;
14'd5901:data <=32'h001CFFD9;14'd5902:data <=32'h0022FFEA;14'd5903:data <=32'h002EFFF4;
14'd5904:data <=32'h003CFFF4;14'd5905:data <=32'h0049FFEE;14'd5906:data <=32'h0052FFE4;
14'd5907:data <=32'h0057FFD5;14'd5908:data <=32'h0057FFC7;14'd5909:data <=32'h0054FFB7;
14'd5910:data <=32'h004FFFA7;14'd5911:data <=32'h0043FF96;14'd5912:data <=32'h0032FF89;
14'd5913:data <=32'h001EFF7F;14'd5914:data <=32'h0005FF7B;14'd5915:data <=32'hFFECFF81;
14'd5916:data <=32'hFFD6FF8C;14'd5917:data <=32'hFFC7FF9F;14'd5918:data <=32'hFFBEFFB4;
14'd5919:data <=32'hFFBEFFC7;14'd5920:data <=32'hFFC2FFD8;14'd5921:data <=32'hFFCBFFE2;
14'd5922:data <=32'hFFD4FFE7;14'd5923:data <=32'hFFDBFFE9;14'd5924:data <=32'hFFDFFFE8;
14'd5925:data <=32'hFFE1FFE8;14'd5926:data <=32'hFFE4FFE9;14'd5927:data <=32'hFFE7FFEB;
14'd5928:data <=32'hFFECFFEB;14'd5929:data <=32'hFFF2FFE9;14'd5930:data <=32'hFFF9FFE4;
14'd5931:data <=32'hFFFCFFDA;14'd5932:data <=32'hFFFDFFCC;14'd5933:data <=32'hFFF9FFBE;
14'd5934:data <=32'hFFEFFFB2;14'd5935:data <=32'hFFE1FFA6;14'd5936:data <=32'hFFCFFF9D;
14'd5937:data <=32'hFFBAFF98;14'd5938:data <=32'hFFA3FF96;14'd5939:data <=32'hFF88FF98;
14'd5940:data <=32'hFF6AFFA0;14'd5941:data <=32'hFF49FFB0;14'd5942:data <=32'hFF2AFFCA;
14'd5943:data <=32'hFF0DFFF1;14'd5944:data <=32'hFEFA0022;14'd5945:data <=32'hFEF5005B;
14'd5946:data <=32'hFF000099;14'd5947:data <=32'hFF1E00D2;14'd5948:data <=32'hFF4A0102;
14'd5949:data <=32'hFF820124;14'd5950:data <=32'hFFC00137;14'd5951:data <=32'hFFFD0139;
14'd5952:data <=32'hFFD10076;14'd5953:data <=32'hFFD60095;14'd5954:data <=32'hFFDD00C2;
14'd5955:data <=32'h001B011E;14'd5956:data <=32'h007E00EC;14'd5957:data <=32'h009E00C6;
14'd5958:data <=32'h00B3009C;14'd5959:data <=32'h00BD0072;14'd5960:data <=32'h00BB0048;
14'd5961:data <=32'h00AF0026;14'd5962:data <=32'h009C000E;14'd5963:data <=32'h00880000;
14'd5964:data <=32'h0078FFF9;14'd5965:data <=32'h006DFFF7;14'd5966:data <=32'h0068FFF7;
14'd5967:data <=32'h0067FFF2;14'd5968:data <=32'h0066FFEB;14'd5969:data <=32'h0062FFE2;
14'd5970:data <=32'h005DFFD9;14'd5971:data <=32'h0053FFD2;14'd5972:data <=32'h004AFFCD;
14'd5973:data <=32'h0041FFCB;14'd5974:data <=32'h003AFFCB;14'd5975:data <=32'h0034FFCB;
14'd5976:data <=32'h0030FFCB;14'd5977:data <=32'h002BFFC9;14'd5978:data <=32'h0026FFC9;
14'd5979:data <=32'h001FFFCA;14'd5980:data <=32'h001AFFCD;14'd5981:data <=32'h0018FFD1;
14'd5982:data <=32'h0019FFD6;14'd5983:data <=32'h001DFFD8;14'd5984:data <=32'h0023FFD6;
14'd5985:data <=32'h0029FFCE;14'd5986:data <=32'h0029FFC3;14'd5987:data <=32'h0025FFB7;
14'd5988:data <=32'h001AFFAC;14'd5989:data <=32'h000BFFA6;14'd5990:data <=32'hFFFAFFA7;
14'd5991:data <=32'hFFECFFAE;14'd5992:data <=32'hFFDFFFBA;14'd5993:data <=32'hFFDCFFC7;
14'd5994:data <=32'hFFDEFFD5;14'd5995:data <=32'hFFE6FFDF;14'd5996:data <=32'hFFF1FFE2;
14'd5997:data <=32'hFFFCFFE2;14'd5998:data <=32'h0006FFDB;14'd5999:data <=32'h000EFFD0;
14'd6000:data <=32'h0012FFC1;14'd6001:data <=32'h0011FFB0;14'd6002:data <=32'h000BFF9C;
14'd6003:data <=32'hFFFFFF86;14'd6004:data <=32'hFFE9FF71;14'd6005:data <=32'hFFCAFF61;
14'd6006:data <=32'hFFA3FF59;14'd6007:data <=32'hFF77FF5D;14'd6008:data <=32'hFF49FF70;
14'd6009:data <=32'hFF1FFF91;14'd6010:data <=32'hFF00FFBF;14'd6011:data <=32'hFEF0FFF4;
14'd6012:data <=32'hFEEF002C;14'd6013:data <=32'hFEFC0061;14'd6014:data <=32'hFF14008E;
14'd6015:data <=32'hFF3400B3;14'd6016:data <=32'hFF36007D;14'd6017:data <=32'hFF3C00AE;
14'd6018:data <=32'hFF4400CF;14'd6019:data <=32'hFF3F00B2;14'd6020:data <=32'hFF9100AD;
14'd6021:data <=32'hFFAA00B8;14'd6022:data <=32'hFFC300BE;14'd6023:data <=32'hFFDD00C1;
14'd6024:data <=32'hFFF400C0;14'd6025:data <=32'h000900BC;14'd6026:data <=32'h001C00B8;
14'd6027:data <=32'h003000B6;14'd6028:data <=32'h004600B4;14'd6029:data <=32'h006000AE;
14'd6030:data <=32'h007C00A2;14'd6031:data <=32'h0099008B;14'd6032:data <=32'h00B0006C;
14'd6033:data <=32'h00BE0047;14'd6034:data <=32'h00C1001F;14'd6035:data <=32'h00B8FFF8;
14'd6036:data <=32'h00A5FFD7;14'd6037:data <=32'h008CFFBF;14'd6038:data <=32'h006FFFAF;
14'd6039:data <=32'h0053FFA8;14'd6040:data <=32'h0038FFA9;14'd6041:data <=32'h0021FFAF;
14'd6042:data <=32'h000DFFB9;14'd6043:data <=32'hFFFDFFCA;14'd6044:data <=32'hFFF2FFDD;
14'd6045:data <=32'hFFF0FFF3;14'd6046:data <=32'hFFF50009;14'd6047:data <=32'h0004001B;
14'd6048:data <=32'h00180026;14'd6049:data <=32'h002F0028;14'd6050:data <=32'h00460020;
14'd6051:data <=32'h0058000F;14'd6052:data <=32'h0062FFFA;14'd6053:data <=32'h0063FFE3;
14'd6054:data <=32'h005DFFD0;14'd6055:data <=32'h0052FFC1;14'd6056:data <=32'h0045FFB8;
14'd6057:data <=32'h0039FFB4;14'd6058:data <=32'h0030FFB2;14'd6059:data <=32'h002AFFB3;
14'd6060:data <=32'h0025FFB2;14'd6061:data <=32'h0022FFAF;14'd6062:data <=32'h001EFFAB;
14'd6063:data <=32'h001BFFA7;14'd6064:data <=32'h0017FFA2;14'd6065:data <=32'h0012FF9D;
14'd6066:data <=32'h000DFF96;14'd6067:data <=32'h0005FF8E;14'd6068:data <=32'hFFFDFF85;
14'd6069:data <=32'hFFEFFF7A;14'd6070:data <=32'hFFDCFF72;14'd6071:data <=32'hFFC4FF6E;
14'd6072:data <=32'hFFA7FF70;14'd6073:data <=32'hFF8CFF7C;14'd6074:data <=32'hFF74FF8F;
14'd6075:data <=32'hFF63FFA8;14'd6076:data <=32'hFF5AFFC4;14'd6077:data <=32'hFF59FFDD;
14'd6078:data <=32'hFF5DFFF2;14'd6079:data <=32'hFF620002;14'd6080:data <=32'hFEF7FFB1;
14'd6081:data <=32'hFED4FFE6;14'd6082:data <=32'hFED40018;14'd6083:data <=32'hFF56FFFB;
14'd6084:data <=32'hFF84FFEE;14'd6085:data <=32'hFF75FFF6;14'd6086:data <=32'hFF690005;
14'd6087:data <=32'hFF5D0019;14'd6088:data <=32'hFF550030;14'd6089:data <=32'hFF50004C;
14'd6090:data <=32'hFF50006D;14'd6091:data <=32'hFF5A0091;14'd6092:data <=32'hFF6D00B7;
14'd6093:data <=32'hFF8C00DA;14'd6094:data <=32'hFFB800F5;14'd6095:data <=32'hFFED0103;
14'd6096:data <=32'h00240100;14'd6097:data <=32'h005800EE;14'd6098:data <=32'h008500CE;
14'd6099:data <=32'h00A400A6;14'd6100:data <=32'h00B60078;14'd6101:data <=32'h00BA004B;
14'd6102:data <=32'h00B40022;14'd6103:data <=32'h00A7FFFE;14'd6104:data <=32'h0092FFE2;
14'd6105:data <=32'h0079FFCA;14'd6106:data <=32'h005EFFBC;14'd6107:data <=32'h003FFFB5;
14'd6108:data <=32'h0022FFB7;14'd6109:data <=32'h0008FFC3;14'd6110:data <=32'hFFF3FFD5;
14'd6111:data <=32'hFFE7FFED;14'd6112:data <=32'hFFE50006;14'd6113:data <=32'hFFEB001C;
14'd6114:data <=32'hFFF8002D;14'd6115:data <=32'h00080037;14'd6116:data <=32'h001A003C;
14'd6117:data <=32'h0029003B;14'd6118:data <=32'h00360039;14'd6119:data <=32'h00430036;
14'd6120:data <=32'h004E0032;14'd6121:data <=32'h005C002E;14'd6122:data <=32'h006B0027;
14'd6123:data <=32'h007C001C;14'd6124:data <=32'h008C000B;14'd6125:data <=32'h0099FFF3;
14'd6126:data <=32'h00A0FFD6;14'd6127:data <=32'h009FFFB7;14'd6128:data <=32'h0097FF99;
14'd6129:data <=32'h0087FF7D;14'd6130:data <=32'h0072FF64;14'd6131:data <=32'h0059FF51;
14'd6132:data <=32'h003CFF41;14'd6133:data <=32'h001DFF38;14'd6134:data <=32'hFFFBFF35;
14'd6135:data <=32'hFFD8FF38;14'd6136:data <=32'hFFB6FF44;14'd6137:data <=32'hFF97FF59;
14'd6138:data <=32'hFF7FFF76;14'd6139:data <=32'hFF72FF98;14'd6140:data <=32'hFF71FFBB;
14'd6141:data <=32'hFF7BFFD8;14'd6142:data <=32'hFF8CFFEC;14'd6143:data <=32'hFFA1FFF6;
14'd6144:data <=32'hFF9CFF48;14'd6145:data <=32'hFF6CFF4B;14'd6146:data <=32'hFF46FF70;
14'd6147:data <=32'hFF8DFFE1;14'd6148:data <=32'hFFC5FFC8;14'd6149:data <=32'hFFBAFFBF;
14'd6150:data <=32'hFFABFFBA;14'd6151:data <=32'hFF99FFB9;14'd6152:data <=32'hFF85FFBE;
14'd6153:data <=32'hFF6FFFC9;14'd6154:data <=32'hFF58FFDB;14'd6155:data <=32'hFF46FFF5;
14'd6156:data <=32'hFF3A0019;14'd6157:data <=32'hFF380042;14'd6158:data <=32'hFF43006B;
14'd6159:data <=32'hFF5C0092;14'd6160:data <=32'hFF7E00AF;14'd6161:data <=32'hFFA500C0;
14'd6162:data <=32'hFFCE00C4;14'd6163:data <=32'hFFF200BE;14'd6164:data <=32'h001200B1;
14'd6165:data <=32'h002A00A0;14'd6166:data <=32'h003D008D;14'd6167:data <=32'h004B007A;
14'd6168:data <=32'h00560067;14'd6169:data <=32'h005C0052;14'd6170:data <=32'h0061003D;
14'd6171:data <=32'h005F0027;14'd6172:data <=32'h00590014;14'd6173:data <=32'h004D0005;
14'd6174:data <=32'h003EFFF9;14'd6175:data <=32'h002EFFF3;14'd6176:data <=32'h0020FFF3;
14'd6177:data <=32'h0015FFF5;14'd6178:data <=32'h000BFFF9;14'd6179:data <=32'h0001FFFE;
14'd6180:data <=32'hFFF80004;14'd6181:data <=32'hFFF0000D;14'd6182:data <=32'hFFE8001B;
14'd6183:data <=32'hFFE3002C;14'd6184:data <=32'hFFE40042;14'd6185:data <=32'hFFEC005B;
14'd6186:data <=32'hFFFF0073;14'd6187:data <=32'h001B0086;14'd6188:data <=32'h00400090;
14'd6189:data <=32'h006A008F;14'd6190:data <=32'h00920081;14'd6191:data <=32'h00B60066;
14'd6192:data <=32'h00D30043;14'd6193:data <=32'h00E50018;14'd6194:data <=32'h00EDFFEB;
14'd6195:data <=32'h00EBFFBD;14'd6196:data <=32'h00DEFF90;14'd6197:data <=32'h00C8FF67;
14'd6198:data <=32'h00A8FF43;14'd6199:data <=32'h0081FF26;14'd6200:data <=32'h0053FF14;
14'd6201:data <=32'h0022FF10;14'd6202:data <=32'hFFF3FF19;14'd6203:data <=32'hFFCBFF2E;
14'd6204:data <=32'hFFAEFF4D;14'd6205:data <=32'hFF9EFF6E;14'd6206:data <=32'hFF9AFF8C;
14'd6207:data <=32'hFFA0FFA4;14'd6208:data <=32'hFFEAFF91;14'd6209:data <=32'hFFE1FF83;
14'd6210:data <=32'hFFC1FF79;14'd6211:data <=32'hFF82FF87;14'd6212:data <=32'hFFB1FF7F;
14'd6213:data <=32'hFFA2FF86;14'd6214:data <=32'hFF94FF90;14'd6215:data <=32'hFF87FF9E;
14'd6216:data <=32'hFF7CFFAD;14'd6217:data <=32'hFF74FFBC;14'd6218:data <=32'hFF6CFFCC;
14'd6219:data <=32'hFF66FFDF;14'd6220:data <=32'hFF62FFF4;14'd6221:data <=32'hFF61000C;
14'd6222:data <=32'hFF690026;14'd6223:data <=32'hFF76003C;14'd6224:data <=32'hFF8B004D;
14'd6225:data <=32'hFFA10056;14'd6226:data <=32'hFFB70057;14'd6227:data <=32'hFFC80051;
14'd6228:data <=32'hFFD20048;14'd6229:data <=32'hFFD50041;14'd6230:data <=32'hFFD4003D;
14'd6231:data <=32'hFFD2003E;14'd6232:data <=32'hFFD20043;14'd6233:data <=32'hFFD6004B;
14'd6234:data <=32'hFFDD0052;14'd6235:data <=32'hFFE70056;14'd6236:data <=32'hFFF20058;
14'd6237:data <=32'hFFFE0057;14'd6238:data <=32'h00090054;14'd6239:data <=32'h0012004E;
14'd6240:data <=32'h001C0047;14'd6241:data <=32'h0023003E;14'd6242:data <=32'h00290032;
14'd6243:data <=32'h002B0024;14'd6244:data <=32'h00270015;14'd6245:data <=32'h001D0007;
14'd6246:data <=32'h000DFFFD;14'd6247:data <=32'hFFF9FFFC;14'd6248:data <=32'hFFE20003;
14'd6249:data <=32'hFFD00015;14'd6250:data <=32'hFFC50030;14'd6251:data <=32'hFFC5004E;
14'd6252:data <=32'hFFD0006D;14'd6253:data <=32'hFFE70088;14'd6254:data <=32'h00040099;
14'd6255:data <=32'h002700A3;14'd6256:data <=32'h004A00A2;14'd6257:data <=32'h006D009A;
14'd6258:data <=32'h008C0089;14'd6259:data <=32'h00A70073;14'd6260:data <=32'h00BE0058;
14'd6261:data <=32'h00CF0038;14'd6262:data <=32'h00DA0014;14'd6263:data <=32'h00DDFFF0;
14'd6264:data <=32'h00D7FFC9;14'd6265:data <=32'h00C9FFA8;14'd6266:data <=32'h00B3FF8C;
14'd6267:data <=32'h009BFF78;14'd6268:data <=32'h0082FF6B;14'd6269:data <=32'h006DFF64;
14'd6270:data <=32'h005DFF5E;14'd6271:data <=32'h004EFF58;14'd6272:data <=32'hFFEFFF7F;
14'd6273:data <=32'hFFEEFF82;14'd6274:data <=32'hFFF4FF79;14'd6275:data <=32'h0031FF1C;
14'd6276:data <=32'h0042FEFD;14'd6277:data <=32'h0011FEF3;14'd6278:data <=32'hFFDEFEF4;
14'd6279:data <=32'hFFADFF03;14'd6280:data <=32'hFF84FF1D;14'd6281:data <=32'hFF61FF3E;
14'd6282:data <=32'hFF48FF62;14'd6283:data <=32'hFF37FF8A;14'd6284:data <=32'hFF2EFFB5;
14'd6285:data <=32'hFF2FFFE0;14'd6286:data <=32'hFF3B000A;14'd6287:data <=32'hFF51002E;
14'd6288:data <=32'hFF71004A;14'd6289:data <=32'hFF960058;14'd6290:data <=32'hFFBB0059;
14'd6291:data <=32'hFFDA004D;14'd6292:data <=32'hFFEF0039;14'd6293:data <=32'hFFF90022;
14'd6294:data <=32'hFFF8000C;14'd6295:data <=32'hFFEEFFFD;14'd6296:data <=32'hFFE1FFF4;
14'd6297:data <=32'hFFD3FFF2;14'd6298:data <=32'hFFC7FFF6;14'd6299:data <=32'hFFBEFFFE;
14'd6300:data <=32'hFFB80008;14'd6301:data <=32'hFFB40013;14'd6302:data <=32'hFFB4001E;
14'd6303:data <=32'hFFB5002A;14'd6304:data <=32'hFFBA0036;14'd6305:data <=32'hFFC30040;
14'd6306:data <=32'hFFD00048;14'd6307:data <=32'hFFDE004A;14'd6308:data <=32'hFFEA0048;
14'd6309:data <=32'hFFF30042;14'd6310:data <=32'hFFF80037;14'd6311:data <=32'hFFF7002F;
14'd6312:data <=32'hFFF00029;14'd6313:data <=32'hFFE70029;14'd6314:data <=32'hFFE0002F;
14'd6315:data <=32'hFFDB003A;14'd6316:data <=32'hFFDB0047;14'd6317:data <=32'hFFE10054;
14'd6318:data <=32'hFFEB005E;14'd6319:data <=32'hFFF80064;14'd6320:data <=32'h00030066;
14'd6321:data <=32'h000D0067;14'd6322:data <=32'h00160066;14'd6323:data <=32'h001E0069;
14'd6324:data <=32'h0026006B;14'd6325:data <=32'h0030006F;14'd6326:data <=32'h003E0071;
14'd6327:data <=32'h004E0072;14'd6328:data <=32'h005F0070;14'd6329:data <=32'h0070006B;
14'd6330:data <=32'h00830063;14'd6331:data <=32'h0094005A;14'd6332:data <=32'h00A9004F;
14'd6333:data <=32'h00BE0040;14'd6334:data <=32'h00D5002A;14'd6335:data <=32'h00EB000B;
14'd6336:data <=32'h0075FF95;14'd6337:data <=32'h0072FF8B;14'd6338:data <=32'h007AFF91;
14'd6339:data <=32'h00EFFFBB;14'd6340:data <=32'h011CFF74;14'd6341:data <=32'h00FBFF3C;
14'd6342:data <=32'h00CEFF0D;14'd6343:data <=32'h0095FEEC;14'd6344:data <=32'h005AFEDC;
14'd6345:data <=32'h0021FED9;14'd6346:data <=32'hFFE9FEE1;14'd6347:data <=32'hFFB6FEF4;
14'd6348:data <=32'hFF88FF13;14'd6349:data <=32'hFF64FF3A;14'd6350:data <=32'hFF4DFF67;
14'd6351:data <=32'hFF42FF99;14'd6352:data <=32'hFF45FFC9;14'd6353:data <=32'hFF55FFF2;
14'd6354:data <=32'hFF700011;14'd6355:data <=32'hFF8E0023;14'd6356:data <=32'hFFAB0029;
14'd6357:data <=32'hFFC20026;14'd6358:data <=32'hFFD3001E;14'd6359:data <=32'hFFDE0014;
14'd6360:data <=32'hFFE3000C;14'd6361:data <=32'hFFE50006;14'd6362:data <=32'hFFE70000;
14'd6363:data <=32'hFFE8FFFB;14'd6364:data <=32'hFFEAFFF5;14'd6365:data <=32'hFFE8FFEE;
14'd6366:data <=32'hFFE4FFE7;14'd6367:data <=32'hFFDCFFE3;14'd6368:data <=32'hFFD2FFE1;
14'd6369:data <=32'hFFC7FFE1;14'd6370:data <=32'hFFBEFFE5;14'd6371:data <=32'hFFB5FFEB;
14'd6372:data <=32'hFFAFFFF4;14'd6373:data <=32'hFFAAFFFB;14'd6374:data <=32'hFFA50003;
14'd6375:data <=32'hFF9F000D;14'd6376:data <=32'hFF990019;14'd6377:data <=32'hFF950029;
14'd6378:data <=32'hFF96003D;14'd6379:data <=32'hFF9B0051;14'd6380:data <=32'hFFA90065;
14'd6381:data <=32'hFFBC0075;14'd6382:data <=32'hFFD4007C;14'd6383:data <=32'hFFEC007C;
14'd6384:data <=32'h00010074;14'd6385:data <=32'h00110067;14'd6386:data <=32'h00170055;
14'd6387:data <=32'h00160047;14'd6388:data <=32'h0010003D;14'd6389:data <=32'h00060039;
14'd6390:data <=32'hFFFC003C;14'd6391:data <=32'hFFF40043;14'd6392:data <=32'hFFF00050;
14'd6393:data <=32'hFFF00060;14'd6394:data <=32'hFFF50073;14'd6395:data <=32'h00000088;
14'd6396:data <=32'h0012009C;14'd6397:data <=32'h002E00AE;14'd6398:data <=32'h005500BA;
14'd6399:data <=32'h008300BB;14'd6400:data <=32'h00850061;14'd6401:data <=32'h00A8005D;
14'd6402:data <=32'h00B60056;14'd6403:data <=32'h00A8007A;14'd6404:data <=32'h00FA0046;
14'd6405:data <=32'h01030015;14'd6406:data <=32'h0100FFE6;14'd6407:data <=32'h00F2FFB9;
14'd6408:data <=32'h00DCFF96;14'd6409:data <=32'h00C2FF76;14'd6410:data <=32'h00A5FF5F;
14'd6411:data <=32'h0086FF4C;14'd6412:data <=32'h0064FF3F;14'd6413:data <=32'h0041FF39;
14'd6414:data <=32'h001DFF3C;14'd6415:data <=32'hFFFFFF46;14'd6416:data <=32'hFFE4FF56;
14'd6417:data <=32'hFFD3FF69;14'd6418:data <=32'hFFC6FF7C;14'd6419:data <=32'hFFC0FF8C;
14'd6420:data <=32'hFFBBFF98;14'd6421:data <=32'hFFB5FFA3;14'd6422:data <=32'hFFAEFFAE;
14'd6423:data <=32'hFFA6FFBA;14'd6424:data <=32'hFFA0FFCC;14'd6425:data <=32'hFF9EFFDF;
14'd6426:data <=32'hFFA3FFF4;14'd6427:data <=32'hFFAF0007;14'd6428:data <=32'hFFC00015;
14'd6429:data <=32'hFFD5001A;14'd6430:data <=32'hFFEA0019;14'd6431:data <=32'hFFFB0010;
14'd6432:data <=32'h00080001;14'd6433:data <=32'h000EFFF1;14'd6434:data <=32'h0010FFDF;
14'd6435:data <=32'h000BFFCE;14'd6436:data <=32'h0001FFBD;14'd6437:data <=32'hFFF3FFAF;
14'd6438:data <=32'hFFDFFFA4;14'd6439:data <=32'hFFC7FF9E;14'd6440:data <=32'hFFABFFA0;
14'd6441:data <=32'hFF8FFFAB;14'd6442:data <=32'hFF75FFBF;14'd6443:data <=32'hFF62FFDA;
14'd6444:data <=32'hFF58FFFC;14'd6445:data <=32'hFF5A001F;14'd6446:data <=32'hFF650040;
14'd6447:data <=32'hFF7A0058;14'd6448:data <=32'hFF920067;14'd6449:data <=32'hFFAA006E;
14'd6450:data <=32'hFFBF006E;14'd6451:data <=32'hFFCE0068;14'd6452:data <=32'hFFD70062;
14'd6453:data <=32'hFFDB005D;14'd6454:data <=32'hFFDD005B;14'd6455:data <=32'hFFDE005C;
14'd6456:data <=32'hFFDF005E;14'd6457:data <=32'hFFE00064;14'd6458:data <=32'hFFE1006B;
14'd6459:data <=32'hFFE40074;14'd6460:data <=32'hFFEA0082;14'd6461:data <=32'hFFF40092;
14'd6462:data <=32'h000600A2;14'd6463:data <=32'h002000AE;14'd6464:data <=32'hFFC300A2;
14'd6465:data <=32'hFFE700D1;14'd6466:data <=32'h001500DE;14'd6467:data <=32'h004F0082;
14'd6468:data <=32'h00990063;14'd6469:data <=32'h009E0045;14'd6470:data <=32'h009A002C;
14'd6471:data <=32'h00900016;14'd6472:data <=32'h0085000A;14'd6473:data <=32'h007C0003;
14'd6474:data <=32'h0078FFFF;14'd6475:data <=32'h0076FFFA;14'd6476:data <=32'h0077FFF4;
14'd6477:data <=32'h0077FFEB;14'd6478:data <=32'h0079FFE2;14'd6479:data <=32'h0078FFD7;
14'd6480:data <=32'h0077FFCC;14'd6481:data <=32'h0076FFC0;14'd6482:data <=32'h0074FFB0;
14'd6483:data <=32'h0070FF9E;14'd6484:data <=32'h0067FF89;14'd6485:data <=32'h0055FF74;
14'd6486:data <=32'h003CFF63;14'd6487:data <=32'h001BFF58;14'd6488:data <=32'hFFF7FF58;
14'd6489:data <=32'hFFD5FF64;14'd6490:data <=32'hFFB8FF7A;14'd6491:data <=32'hFFA5FF99;
14'd6492:data <=32'hFF9CFFB9;14'd6493:data <=32'hFF9FFFD9;14'd6494:data <=32'hFFACFFF2;
14'd6495:data <=32'hFFBD0005;14'd6496:data <=32'hFFD20010;14'd6497:data <=32'hFFE60015;
14'd6498:data <=32'hFFFB0013;14'd6499:data <=32'h000D000B;14'd6500:data <=32'h001DFFFD;
14'd6501:data <=32'h0028FFEB;14'd6502:data <=32'h002DFFD5;14'd6503:data <=32'h002AFFBD;
14'd6504:data <=32'h001FFFA5;14'd6505:data <=32'h000DFF92;14'd6506:data <=32'hFFF4FF85;
14'd6507:data <=32'hFFD8FF80;14'd6508:data <=32'hFFBDFF84;14'd6509:data <=32'hFFA6FF8F;
14'd6510:data <=32'hFF92FF9F;14'd6511:data <=32'hFF84FFB0;14'd6512:data <=32'hFF7CFFBF;
14'd6513:data <=32'hFF74FFCD;14'd6514:data <=32'hFF6CFFDA;14'd6515:data <=32'hFF63FFE8;
14'd6516:data <=32'hFF58FFF9;14'd6517:data <=32'hFF4F000F;14'd6518:data <=32'hFF4A0029;
14'd6519:data <=32'hFF4A0048;14'd6520:data <=32'hFF500066;14'd6521:data <=32'hFF5F0083;
14'd6522:data <=32'hFF73009D;14'd6523:data <=32'hFF8B00B2;14'd6524:data <=32'hFFA600C4;
14'd6525:data <=32'hFFC400D1;14'd6526:data <=32'hFFE500DA;14'd6527:data <=32'h000900DC;
14'd6528:data <=32'hFF7A0032;14'd6529:data <=32'hFF71006D;14'd6530:data <=32'hFF8F00A7;
14'd6531:data <=32'h003F00C3;14'd6532:data <=32'h0094009A;14'd6533:data <=32'h009D006E;
14'd6534:data <=32'h00980045;14'd6535:data <=32'h00890023;14'd6536:data <=32'h0072000F;
14'd6537:data <=32'h005A0005;14'd6538:data <=32'h00470005;14'd6539:data <=32'h0039000D;
14'd6540:data <=32'h00320016;14'd6541:data <=32'h00310021;14'd6542:data <=32'h00350029;
14'd6543:data <=32'h003D0031;14'd6544:data <=32'h00490035;14'd6545:data <=32'h00580036;
14'd6546:data <=32'h006C0031;14'd6547:data <=32'h007E0025;14'd6548:data <=32'h008F0010;
14'd6549:data <=32'h0099FFF4;14'd6550:data <=32'h009AFFD3;14'd6551:data <=32'h0090FFB4;
14'd6552:data <=32'h007BFF99;14'd6553:data <=32'h005FFF86;14'd6554:data <=32'h0040FF7E;
14'd6555:data <=32'h0024FF80;14'd6556:data <=32'h000CFF89;14'd6557:data <=32'hFFF9FF96;
14'd6558:data <=32'hFFEDFFA5;14'd6559:data <=32'hFFE6FFB3;14'd6560:data <=32'hFFE3FFC1;
14'd6561:data <=32'hFFE2FFCE;14'd6562:data <=32'hFFE2FFD9;14'd6563:data <=32'hFFE6FFE4;
14'd6564:data <=32'hFFEDFFEE;14'd6565:data <=32'hFFF7FFF4;14'd6566:data <=32'h0004FFF8;
14'd6567:data <=32'h0010FFF8;14'd6568:data <=32'h001CFFF0;14'd6569:data <=32'h0024FFE7;
14'd6570:data <=32'h002BFFDB;14'd6571:data <=32'h002DFFCC;14'd6572:data <=32'h002CFFC0;
14'd6573:data <=32'h002AFFB2;14'd6574:data <=32'h0027FFA5;14'd6575:data <=32'h0022FF95;
14'd6576:data <=32'h0019FF83;14'd6577:data <=32'h000BFF6D;14'd6578:data <=32'hFFF4FF59;
14'd6579:data <=32'hFFD4FF47;14'd6580:data <=32'hFFAAFF3E;14'd6581:data <=32'hFF7CFF41;
14'd6582:data <=32'hFF4CFF53;14'd6583:data <=32'hFF20FF71;14'd6584:data <=32'hFEFEFF9B;
14'd6585:data <=32'hFEE7FFD0;14'd6586:data <=32'hFEDC0007;14'd6587:data <=32'hFEDE003E;
14'd6588:data <=32'hFEED0074;14'd6589:data <=32'hFF0600A7;14'd6590:data <=32'hFF2B00D3;
14'd6591:data <=32'hFF5800F7;14'd6592:data <=32'hFF830028;14'd6593:data <=32'hFF70004C;
14'd6594:data <=32'hFF640081;14'd6595:data <=32'hFF8B00FD;14'd6596:data <=32'hFFFA00F3;
14'd6597:data <=32'h002200DA;14'd6598:data <=32'h003E00BC;14'd6599:data <=32'h004E009C;
14'd6600:data <=32'h00520080;14'd6601:data <=32'h0051006A;14'd6602:data <=32'h004D005B;
14'd6603:data <=32'h004A0051;14'd6604:data <=32'h0049004A;14'd6605:data <=32'h00470044;
14'd6606:data <=32'h0047003E;14'd6607:data <=32'h00480039;14'd6608:data <=32'h00470035;
14'd6609:data <=32'h00470033;14'd6610:data <=32'h004B0032;14'd6611:data <=32'h0050002F;
14'd6612:data <=32'h00590029;14'd6613:data <=32'h0061001F;14'd6614:data <=32'h00650012;
14'd6615:data <=32'h00640002;14'd6616:data <=32'h005FFFF4;14'd6617:data <=32'h0055FFE9;
14'd6618:data <=32'h0049FFE4;14'd6619:data <=32'h0040FFE3;14'd6620:data <=32'h0039FFE7;
14'd6621:data <=32'h0038FFEA;14'd6622:data <=32'h003AFFEB;14'd6623:data <=32'h003EFFE9;
14'd6624:data <=32'h0041FFE3;14'd6625:data <=32'h0040FFDA;14'd6626:data <=32'h003CFFCF;
14'd6627:data <=32'h0034FFC8;14'd6628:data <=32'h0029FFC4;14'd6629:data <=32'h001FFFC4;
14'd6630:data <=32'h0016FFC7;14'd6631:data <=32'h000FFFCD;14'd6632:data <=32'h000BFFD3;
14'd6633:data <=32'h0009FFDB;14'd6634:data <=32'h000AFFE2;14'd6635:data <=32'h000EFFEA;
14'd6636:data <=32'h0015FFF1;14'd6637:data <=32'h0022FFF4;14'd6638:data <=32'h0031FFF4;
14'd6639:data <=32'h0044FFEF;14'd6640:data <=32'h0057FFDE;14'd6641:data <=32'h0067FFC5;
14'd6642:data <=32'h006FFFA3;14'd6643:data <=32'h006AFF7B;14'd6644:data <=32'h0057FF53;
14'd6645:data <=32'h0036FF2F;14'd6646:data <=32'h000AFF17;14'd6647:data <=32'hFFD7FF0B;
14'd6648:data <=32'hFFA2FF0D;14'd6649:data <=32'hFF6FFF1E;14'd6650:data <=32'hFF42FF39;
14'd6651:data <=32'hFF1EFF5E;14'd6652:data <=32'hFF01FF88;14'd6653:data <=32'hFEEDFFB9;
14'd6654:data <=32'hFEE4FFEC;14'd6655:data <=32'hFEE6001F;14'd6656:data <=32'hFF1AFFF7;
14'd6657:data <=32'hFF060024;14'd6658:data <=32'hFEFA0045;14'd6659:data <=32'hFEF40039;
14'd6660:data <=32'hFF430057;14'd6661:data <=32'hFF560067;14'd6662:data <=32'hFF670074;
14'd6663:data <=32'hFF76007F;14'd6664:data <=32'hFF830089;14'd6665:data <=32'hFF8F0099;
14'd6666:data <=32'hFFA100AA;14'd6667:data <=32'hFFB700B9;14'd6668:data <=32'hFFD400C6;
14'd6669:data <=32'hFFF600C9;14'd6670:data <=32'h001900C5;14'd6671:data <=32'h003700B7;
14'd6672:data <=32'h005300A4;14'd6673:data <=32'h0067008D;14'd6674:data <=32'h00750073;
14'd6675:data <=32'h007F005A;14'd6676:data <=32'h0082003F;14'd6677:data <=32'h00810024;
14'd6678:data <=32'h0079000A;14'd6679:data <=32'h006BFFF3;14'd6680:data <=32'h0056FFE1;
14'd6681:data <=32'h003DFFD9;14'd6682:data <=32'h0023FFDA;14'd6683:data <=32'h000DFFE4;
14'd6684:data <=32'hFFFDFFF7;14'd6685:data <=32'hFFF9000D;14'd6686:data <=32'hFFFE0021;
14'd6687:data <=32'h000B0031;14'd6688:data <=32'h001D003A;14'd6689:data <=32'h0030003A;
14'd6690:data <=32'h00400034;14'd6691:data <=32'h004C0029;14'd6692:data <=32'h0054001C;
14'd6693:data <=32'h0058000F;14'd6694:data <=32'h00580003;14'd6695:data <=32'h0058FFF8;
14'd6696:data <=32'h0054FFEE;14'd6697:data <=32'h004FFFE7;14'd6698:data <=32'h004AFFE0;
14'd6699:data <=32'h0043FFDC;14'd6700:data <=32'h003EFFDC;14'd6701:data <=32'h0039FFDE;
14'd6702:data <=32'h0039FFE2;14'd6703:data <=32'h003FFFE6;14'd6704:data <=32'h0049FFE6;
14'd6705:data <=32'h0056FFDF;14'd6706:data <=32'h0062FFD1;14'd6707:data <=32'h006AFFBB;
14'd6708:data <=32'h006AFFA1;14'd6709:data <=32'h0061FF86;14'd6710:data <=32'h004FFF6D;
14'd6711:data <=32'h0036FF5A;14'd6712:data <=32'h001AFF50;14'd6713:data <=32'hFFFEFF4C;
14'd6714:data <=32'hFFE4FF4E;14'd6715:data <=32'hFFCCFF54;14'd6716:data <=32'hFFB6FF5B;
14'd6717:data <=32'hFFA3FF64;14'd6718:data <=32'hFF90FF70;14'd6719:data <=32'hFF7DFF7F;
14'd6720:data <=32'hFF3AFF2F;14'd6721:data <=32'hFF05FF50;14'd6722:data <=32'hFEF0FF7B;
14'd6723:data <=32'hFF6BFF85;14'd6724:data <=32'hFF99FF8D;14'd6725:data <=32'hFF86FF8E;
14'd6726:data <=32'hFF6EFF92;14'd6727:data <=32'hFF54FF9D;14'd6728:data <=32'hFF36FFB1;
14'd6729:data <=32'hFF1AFFD2;14'd6730:data <=32'hFF07FFFD;14'd6731:data <=32'hFF010030;
14'd6732:data <=32'hFF0A0065;14'd6733:data <=32'hFF220096;14'd6734:data <=32'hFF4700BE;
14'd6735:data <=32'hFF7400DA;14'd6736:data <=32'hFFA400EA;14'd6737:data <=32'hFFD500EE;
14'd6738:data <=32'h000300E7;14'd6739:data <=32'h002D00D6;14'd6740:data <=32'h005200BE;
14'd6741:data <=32'h006F009D;14'd6742:data <=32'h00840077;14'd6743:data <=32'h008B004E;
14'd6744:data <=32'h00880026;14'd6745:data <=32'h00770002;14'd6746:data <=32'h005EFFE7;
14'd6747:data <=32'h003EFFD9;14'd6748:data <=32'h0020FFD7;14'd6749:data <=32'h0005FFDE;
14'd6750:data <=32'hFFF2FFEE;14'd6751:data <=32'hFFE70001;14'd6752:data <=32'hFFE40013;
14'd6753:data <=32'hFFE60023;14'd6754:data <=32'hFFEC0030;14'd6755:data <=32'hFFF2003A;
14'd6756:data <=32'hFFF90043;14'd6757:data <=32'h0002004C;14'd6758:data <=32'h000E0055;
14'd6759:data <=32'h001C005B;14'd6760:data <=32'h002C005F;14'd6761:data <=32'h003E005F;
14'd6762:data <=32'h0052005B;14'd6763:data <=32'h00630052;14'd6764:data <=32'h00730046;
14'd6765:data <=32'h007F0038;14'd6766:data <=32'h008B0028;14'd6767:data <=32'h00950017;
14'd6768:data <=32'h009C0004;14'd6769:data <=32'h00A3FFEE;14'd6770:data <=32'h00A6FFD4;
14'd6771:data <=32'h00A3FFB6;14'd6772:data <=32'h0099FF99;14'd6773:data <=32'h0084FF7E;
14'd6774:data <=32'h0069FF68;14'd6775:data <=32'h0049FF5D;14'd6776:data <=32'h0028FF5B;
14'd6777:data <=32'h000BFF65;14'd6778:data <=32'hFFF6FF74;14'd6779:data <=32'hFFEAFF85;
14'd6780:data <=32'hFFE5FF95;14'd6781:data <=32'hFFE6FFA2;14'd6782:data <=32'hFFEAFFA9;
14'd6783:data <=32'hFFEFFFAB;14'd6784:data <=32'h0013FF13;14'd6785:data <=32'hFFE2FF02;
14'd6786:data <=32'hFFB1FF17;14'd6787:data <=32'hFFD7FF9A;14'd6788:data <=32'h0014FF94;
14'd6789:data <=32'h000DFF7F;14'd6790:data <=32'hFFFDFF68;14'd6791:data <=32'hFFE3FF55;
14'd6792:data <=32'hFFBEFF49;14'd6793:data <=32'hFF94FF49;14'd6794:data <=32'hFF67FF59;
14'd6795:data <=32'hFF40FF76;14'd6796:data <=32'hFF23FF9F;14'd6797:data <=32'hFF14FFCD;
14'd6798:data <=32'hFF11FFFD;14'd6799:data <=32'hFF1A0029;14'd6800:data <=32'hFF2B004F;
14'd6801:data <=32'hFF44006F;14'd6802:data <=32'hFF610088;14'd6803:data <=32'hFF80009B;
14'd6804:data <=32'hFFA300A7;14'd6805:data <=32'hFFC600AB;14'd6806:data <=32'hFFE900A7;
14'd6807:data <=32'h0008009A;14'd6808:data <=32'h00220086;14'd6809:data <=32'h0032006E;
14'd6810:data <=32'h003B0055;14'd6811:data <=32'h003B003D;14'd6812:data <=32'h0035002B;
14'd6813:data <=32'h002D001D;14'd6814:data <=32'h00250014;14'd6815:data <=32'h001D000D;
14'd6816:data <=32'h00160008;14'd6817:data <=32'h000E0001;14'd6818:data <=32'h0004FFFB;
14'd6819:data <=32'hFFF6FFF8;14'd6820:data <=32'hFFE5FFF9;14'd6821:data <=32'hFFD20001;
14'd6822:data <=32'hFFC30011;14'd6823:data <=32'hFFB70028;14'd6824:data <=32'hFFB40043;
14'd6825:data <=32'hFFB9005F;14'd6826:data <=32'hFFC7007A;14'd6827:data <=32'hFFDD0093;
14'd6828:data <=32'hFFF900A5;14'd6829:data <=32'h001A00B1;14'd6830:data <=32'h003E00B4;
14'd6831:data <=32'h006300B1;14'd6832:data <=32'h008900A5;14'd6833:data <=32'h00AE008F;
14'd6834:data <=32'h00CE006F;14'd6835:data <=32'h00E70045;14'd6836:data <=32'h00F40016;
14'd6837:data <=32'h00F3FFE3;14'd6838:data <=32'h00E2FFB3;14'd6839:data <=32'h00C7FF8C;
14'd6840:data <=32'h00A2FF6F;14'd6841:data <=32'h007AFF61;14'd6842:data <=32'h0056FF5F;
14'd6843:data <=32'h0037FF67;14'd6844:data <=32'h0020FF75;14'd6845:data <=32'h0012FF84;
14'd6846:data <=32'h000AFF92;14'd6847:data <=32'h0007FF9C;14'd6848:data <=32'h004DFF9E;
14'd6849:data <=32'h004BFF89;14'd6850:data <=32'h0031FF74;14'd6851:data <=32'hFFEEFF7A;
14'd6852:data <=32'h0023FF82;14'd6853:data <=32'h001DFF7B;14'd6854:data <=32'h0014FF71;
14'd6855:data <=32'h0005FF68;14'd6856:data <=32'hFFF0FF5E;14'd6857:data <=32'hFFD6FF5B;
14'd6858:data <=32'hFFB8FF60;14'd6859:data <=32'hFF9DFF6E;14'd6860:data <=32'hFF87FF85;
14'd6861:data <=32'hFF79FF9F;14'd6862:data <=32'hFF74FFBA;14'd6863:data <=32'hFF77FFD1;
14'd6864:data <=32'hFF7CFFE3;14'd6865:data <=32'hFF83FFF1;14'd6866:data <=32'hFF8AFFFB;
14'd6867:data <=32'hFF8E0004;14'd6868:data <=32'hFF91000E;14'd6869:data <=32'hFF960018;
14'd6870:data <=32'hFF9C0021;14'd6871:data <=32'hFFA40029;14'd6872:data <=32'hFFAB002F;
14'd6873:data <=32'hFFB20034;14'd6874:data <=32'hFFB90038;14'd6875:data <=32'hFFBF003C;
14'd6876:data <=32'hFFC50042;14'd6877:data <=32'hFFCE0048;14'd6878:data <=32'hFFDA0050;
14'd6879:data <=32'hFFE90051;14'd6880:data <=32'hFFFA004F;14'd6881:data <=32'h000C0045;
14'd6882:data <=32'h00180034;14'd6883:data <=32'h001D001F;14'd6884:data <=32'h00190007;
14'd6885:data <=32'h000BFFF4;14'd6886:data <=32'hFFF6FFE9;14'd6887:data <=32'hFFDCFFE6;
14'd6888:data <=32'hFFC2FFED;14'd6889:data <=32'hFFACFFFD;14'd6890:data <=32'hFF9C0014;
14'd6891:data <=32'hFF93002F;14'd6892:data <=32'hFF92004D;14'd6893:data <=32'hFF98006D;
14'd6894:data <=32'hFFA6008A;14'd6895:data <=32'hFFBC00A6;14'd6896:data <=32'hFFD900BD;
14'd6897:data <=32'hFFFE00CD;14'd6898:data <=32'h002700D3;14'd6899:data <=32'h005200CF;
14'd6900:data <=32'h007B00BE;14'd6901:data <=32'h009D00A4;14'd6902:data <=32'h00B60082;
14'd6903:data <=32'h00C4005D;14'd6904:data <=32'h00C8003A;14'd6905:data <=32'h00C4001C;
14'd6906:data <=32'h00BD0005;14'd6907:data <=32'h00B6FFF2;14'd6908:data <=32'h00B0FFE2;
14'd6909:data <=32'h00ACFFD2;14'd6910:data <=32'h00A8FFC0;14'd6911:data <=32'h00A2FFAD;
14'd6912:data <=32'h0035FFB2;14'd6913:data <=32'h0037FFB7;14'd6914:data <=32'h0043FFAF;
14'd6915:data <=32'h0093FF6B;14'd6916:data <=32'h00B5FF5C;14'd6917:data <=32'h0098FF41;
14'd6918:data <=32'h0075FF2A;14'd6919:data <=32'h0050FF1B;14'd6920:data <=32'h0025FF14;
14'd6921:data <=32'hFFF9FF15;14'd6922:data <=32'hFFCDFF23;14'd6923:data <=32'hFFA6FF3C;
14'd6924:data <=32'hFF88FF5F;14'd6925:data <=32'hFF78FF88;14'd6926:data <=32'hFF75FFB0;
14'd6927:data <=32'hFF7FFFD3;14'd6928:data <=32'hFF93FFEE;14'd6929:data <=32'hFFA9FFFC;
14'd6930:data <=32'hFFBF0001;14'd6931:data <=32'hFFD0FFFE;14'd6932:data <=32'hFFDCFFF7;
14'd6933:data <=32'hFFE2FFEE;14'd6934:data <=32'hFFE5FFE5;14'd6935:data <=32'hFFE3FFDC;
14'd6936:data <=32'hFFDEFFD4;14'd6937:data <=32'hFFD4FFCF;14'd6938:data <=32'hFFC8FFCC;
14'd6939:data <=32'hFFBAFFCE;14'd6940:data <=32'hFFABFFD6;14'd6941:data <=32'hFF9EFFE4;
14'd6942:data <=32'hFF98FFF8;14'd6943:data <=32'hFF99000D;14'd6944:data <=32'hFFA10020;
14'd6945:data <=32'hFFB0002E;14'd6946:data <=32'hFFC30034;14'd6947:data <=32'hFFD40032;
14'd6948:data <=32'hFFE2002A;14'd6949:data <=32'hFFE8001F;14'd6950:data <=32'hFFE90012;
14'd6951:data <=32'hFFE3000A;14'd6952:data <=32'hFFDB0005;14'd6953:data <=32'hFFD00003;
14'd6954:data <=32'hFFC60007;14'd6955:data <=32'hFFBE000C;14'd6956:data <=32'hFFB80014;
14'd6957:data <=32'hFFB2001D;14'd6958:data <=32'hFFAD0028;14'd6959:data <=32'hFFA90035;
14'd6960:data <=32'hFFA80045;14'd6961:data <=32'hFFAA0056;14'd6962:data <=32'hFFB10067;
14'd6963:data <=32'hFFBD0078;14'd6964:data <=32'hFFCC0085;14'd6965:data <=32'hFFDC008E;
14'd6966:data <=32'hFFED0094;14'd6967:data <=32'hFFFB0099;14'd6968:data <=32'h000800A0;
14'd6969:data <=32'h001700A7;14'd6970:data <=32'h002A00B0;14'd6971:data <=32'h004400BA;
14'd6972:data <=32'h006400BE;14'd6973:data <=32'h008A00BB;14'd6974:data <=32'h00B400AC;
14'd6975:data <=32'h00DB0092;14'd6976:data <=32'h0083FFE9;14'd6977:data <=32'h0082FFE5;
14'd6978:data <=32'h0087FFF5;14'd6979:data <=32'h00F30044;14'd6980:data <=32'h013A001C;
14'd6981:data <=32'h013AFFE0;14'd6982:data <=32'h012CFFA5;14'd6983:data <=32'h0112FF6E;
14'd6984:data <=32'h00EBFF3E;14'd6985:data <=32'h00B9FF18;14'd6986:data <=32'h007FFF01;
14'd6987:data <=32'h0042FEFA;14'd6988:data <=32'h0008FF06;14'd6989:data <=32'hFFD8FF20;
14'd6990:data <=32'hFFB5FF46;14'd6991:data <=32'hFFA0FF6D;14'd6992:data <=32'hFF9BFF93;
14'd6993:data <=32'hFF9EFFB4;14'd6994:data <=32'hFFAAFFCC;14'd6995:data <=32'hFFB7FFDD;
14'd6996:data <=32'hFFC4FFE8;14'd6997:data <=32'hFFD2FFEF;14'd6998:data <=32'hFFDDFFF1;
14'd6999:data <=32'hFFE8FFF1;14'd7000:data <=32'hFFF2FFEE;14'd7001:data <=32'hFFFAFFE7;
14'd7002:data <=32'hFFFEFFDC;14'd7003:data <=32'hFFFDFFD2;14'd7004:data <=32'hFFF6FFC9;
14'd7005:data <=32'hFFEDFFC3;14'd7006:data <=32'hFFE1FFC2;14'd7007:data <=32'hFFD8FFC5;
14'd7008:data <=32'hFFD1FFCB;14'd7009:data <=32'hFFCEFFD0;14'd7010:data <=32'hFFCCFFD3;
14'd7011:data <=32'hFFCBFFD4;14'd7012:data <=32'hFFC8FFD3;14'd7013:data <=32'hFFC2FFD2;
14'd7014:data <=32'hFFB6FFD2;14'd7015:data <=32'hFFABFFD7;14'd7016:data <=32'hFF9FFFE2;
14'd7017:data <=32'hFF97FFF0;14'd7018:data <=32'hFF940002;14'd7019:data <=32'hFF960013;
14'd7020:data <=32'hFF9E0023;14'd7021:data <=32'hFFA9002D;14'd7022:data <=32'hFFB50032;
14'd7023:data <=32'hFFBF0033;14'd7024:data <=32'hFFC70031;14'd7025:data <=32'hFFCC002E;
14'd7026:data <=32'hFFCF002B;14'd7027:data <=32'hFFCF0027;14'd7028:data <=32'hFFCB0024;
14'd7029:data <=32'hFFC40021;14'd7030:data <=32'hFFBA0021;14'd7031:data <=32'hFFAC0026;
14'd7032:data <=32'hFF9C0032;14'd7033:data <=32'hFF8D0048;14'd7034:data <=32'hFF840068;
14'd7035:data <=32'hFF85008F;14'd7036:data <=32'hFF9400BA;14'd7037:data <=32'hFFB300E1;
14'd7038:data <=32'hFFDF0100;14'd7039:data <=32'h00150113;14'd7040:data <=32'h00410098;
14'd7041:data <=32'h005B00A3;14'd7042:data <=32'h006100A9;14'd7043:data <=32'h004900DC;
14'd7044:data <=32'h00AE00D6;14'd7045:data <=32'h00D100B4;14'd7046:data <=32'h00EC008A;
14'd7047:data <=32'h0100005D;14'd7048:data <=32'h0108002C;14'd7049:data <=32'h0104FFFA;
14'd7050:data <=32'h00F4FFCC;14'd7051:data <=32'h00DBFFA4;14'd7052:data <=32'h00B9FF89;
14'd7053:data <=32'h0096FF78;14'd7054:data <=32'h0076FF73;14'd7055:data <=32'h005AFF74;
14'd7056:data <=32'h0044FF77;14'd7057:data <=32'h0034FF7B;14'd7058:data <=32'h0025FF7E;
14'd7059:data <=32'h0017FF80;14'd7060:data <=32'h0007FF83;14'd7061:data <=32'hFFF6FF89;
14'd7062:data <=32'hFFE6FF94;14'd7063:data <=32'hFFD9FFA2;14'd7064:data <=32'hFFD1FFB3;
14'd7065:data <=32'hFFCFFFC5;14'd7066:data <=32'hFFD1FFD4;14'd7067:data <=32'hFFD6FFE0;
14'd7068:data <=32'hFFDFFFEA;14'd7069:data <=32'hFFE7FFF1;14'd7070:data <=32'hFFF0FFF6;
14'd7071:data <=32'hFFFCFFF8;14'd7072:data <=32'h0008FFF7;14'd7073:data <=32'h0015FFF1;
14'd7074:data <=32'h0021FFE6;14'd7075:data <=32'h0029FFD4;14'd7076:data <=32'h002BFFBE;
14'd7077:data <=32'h0023FFA6;14'd7078:data <=32'h0012FF91;14'd7079:data <=32'hFFF9FF82;
14'd7080:data <=32'hFFDCFF7C;14'd7081:data <=32'hFFBDFF81;14'd7082:data <=32'hFFA1FF8E;
14'd7083:data <=32'hFF8DFFA4;14'd7084:data <=32'hFF80FFBD;14'd7085:data <=32'hFF7BFFD5;
14'd7086:data <=32'hFF7DFFEC;14'd7087:data <=32'hFF83FFFE;14'd7088:data <=32'hFF8C000C;
14'd7089:data <=32'hFF960017;14'd7090:data <=32'hFF9F001E;14'd7091:data <=32'hFFAA0020;
14'd7092:data <=32'hFFB20021;14'd7093:data <=32'hFFB8001C;14'd7094:data <=32'hFFB90017;
14'd7095:data <=32'hFFB30011;14'd7096:data <=32'hFFA9000D;14'd7097:data <=32'hFF980010;
14'd7098:data <=32'hFF85001E;14'd7099:data <=32'hFF760034;14'd7100:data <=32'hFF6D0055;
14'd7101:data <=32'hFF710078;14'd7102:data <=32'hFF81009C;14'd7103:data <=32'hFF9B00BB;
14'd7104:data <=32'hFF690084;14'd7105:data <=32'hFF7500BA;14'd7106:data <=32'hFF9000D5;
14'd7107:data <=32'hFFD1009C;14'd7108:data <=32'h001F00AB;14'd7109:data <=32'h003100A1;
14'd7110:data <=32'h00420096;14'd7111:data <=32'h004E008B;14'd7112:data <=32'h005C007F;
14'd7113:data <=32'h00660071;14'd7114:data <=32'h006E0063;14'd7115:data <=32'h00730055;
14'd7116:data <=32'h00740049;14'd7117:data <=32'h00780041;14'd7118:data <=32'h007C003B;
14'd7119:data <=32'h00860035;14'd7120:data <=32'h0093002B;14'd7121:data <=32'h00A1001A;
14'd7122:data <=32'h00AC0001;14'd7123:data <=32'h00B0FFE2;14'd7124:data <=32'h00AAFFC0;
14'd7125:data <=32'h0099FFA0;14'd7126:data <=32'h0080FF87;14'd7127:data <=32'h0060FF76;
14'd7128:data <=32'h003FFF70;14'd7129:data <=32'h001FFF72;14'd7130:data <=32'h0003FF7B;
14'd7131:data <=32'hFFEBFF8A;14'd7132:data <=32'hFFDAFF9F;14'd7133:data <=32'hFFCDFFB6;
14'd7134:data <=32'hFFC8FFCF;14'd7135:data <=32'hFFCAFFE8;14'd7136:data <=32'hFFD4FFFF;
14'd7137:data <=32'hFFE70012;14'd7138:data <=32'h0000001D;14'd7139:data <=32'h001B001D;
14'd7140:data <=32'h00350014;14'd7141:data <=32'h004A0000;14'd7142:data <=32'h0056FFE6;
14'd7143:data <=32'h0058FFC9;14'd7144:data <=32'h0050FFAE;14'd7145:data <=32'h0041FF98;
14'd7146:data <=32'h002EFF88;14'd7147:data <=32'h0019FF7D;14'd7148:data <=32'h0004FF7A;
14'd7149:data <=32'hFFF2FF79;14'd7150:data <=32'hFFE0FF7B;14'd7151:data <=32'hFFD0FF7C;
14'd7152:data <=32'hFFBFFF7F;14'd7153:data <=32'hFFADFF83;14'd7154:data <=32'hFF9CFF8C;
14'd7155:data <=32'hFF8BFF97;14'd7156:data <=32'hFF7BFFA4;14'd7157:data <=32'hFF6FFFB4;
14'd7158:data <=32'hFF66FFC4;14'd7159:data <=32'hFF5CFFD6;14'd7160:data <=32'hFF54FFE7;
14'd7161:data <=32'hFF4CFFFC;14'd7162:data <=32'hFF450014;14'd7163:data <=32'hFF42002F;
14'd7164:data <=32'hFF450050;14'd7165:data <=32'hFF510072;14'd7166:data <=32'hFF680090;
14'd7167:data <=32'hFF8600A7;14'd7168:data <=32'hFF50FFDC;14'd7169:data <=32'hFF2B000B;
14'd7170:data <=32'hFF290047;14'd7171:data <=32'hFFBE0098;14'd7172:data <=32'h000E009E;
14'd7173:data <=32'h001E0085;14'd7174:data <=32'h0025006F;14'd7175:data <=32'h0024005C;
14'd7176:data <=32'h0020004E;14'd7177:data <=32'h001A0045;14'd7178:data <=32'h0011003E;
14'd7179:data <=32'h0007003F;14'd7180:data <=32'hFFFE0045;14'd7181:data <=32'hFFF90052;
14'd7182:data <=32'hFFFA0063;14'd7183:data <=32'h00050077;14'd7184:data <=32'h001A0088;
14'd7185:data <=32'h00380091;14'd7186:data <=32'h005A008E;14'd7187:data <=32'h007C0080;
14'd7188:data <=32'h00980066;14'd7189:data <=32'h00AA0044;14'd7190:data <=32'h00B10020;
14'd7191:data <=32'h00ADFFFD;14'd7192:data <=32'h00A1FFDF;14'd7193:data <=32'h0090FFC6;
14'd7194:data <=32'h007BFFB4;14'd7195:data <=32'h0063FFA6;14'd7196:data <=32'h004BFF9F;
14'd7197:data <=32'h0032FF9D;14'd7198:data <=32'h001CFFA1;14'd7199:data <=32'h0007FFAC;
14'd7200:data <=32'hFFF6FFBC;14'd7201:data <=32'hFFECFFD0;14'd7202:data <=32'hFFEBFFE5;
14'd7203:data <=32'hFFF1FFF8;14'd7204:data <=32'hFFFD0006;14'd7205:data <=32'h000B000F;
14'd7206:data <=32'h001B0010;14'd7207:data <=32'h0029000D;14'd7208:data <=32'h00340007;
14'd7209:data <=32'h003D0001;14'd7210:data <=32'h0045FFFB;14'd7211:data <=32'h004EFFF3;
14'd7212:data <=32'h0057FFEA;14'd7213:data <=32'h0063FFDC;14'd7214:data <=32'h006CFFC8;
14'd7215:data <=32'h0073FFAF;14'd7216:data <=32'h0073FF90;14'd7217:data <=32'h0068FF70;
14'd7218:data <=32'h0054FF50;14'd7219:data <=32'h0037FF34;14'd7220:data <=32'h0012FF20;
14'd7221:data <=32'hFFE9FF15;14'd7222:data <=32'hFFBDFF13;14'd7223:data <=32'hFF8FFF1A;
14'd7224:data <=32'hFF63FF29;14'd7225:data <=32'hFF39FF42;14'd7226:data <=32'hFF13FF66;
14'd7227:data <=32'hFEF3FF94;14'd7228:data <=32'hFEE0FFCC;14'd7229:data <=32'hFEDD0007;
14'd7230:data <=32'hFEE80042;14'd7231:data <=32'hFF050077;14'd7232:data <=32'hFF86FFC4;
14'd7233:data <=32'hFF63FFD3;14'd7234:data <=32'hFF3DFFF6;14'd7235:data <=32'hFF330080;
14'd7236:data <=32'hFF8F00A1;14'd7237:data <=32'hFFB0009C;14'd7238:data <=32'hFFCA0092;
14'd7239:data <=32'hFFDC0085;14'd7240:data <=32'hFFEC0079;14'd7241:data <=32'hFFF5006C;
14'd7242:data <=32'hFFFB0060;14'd7243:data <=32'hFFFB0054;14'd7244:data <=32'hFFF7004C;
14'd7245:data <=32'hFFF1004A;14'd7246:data <=32'hFFEB004E;14'd7247:data <=32'hFFE80058;
14'd7248:data <=32'hFFED0066;14'd7249:data <=32'hFFF90073;14'd7250:data <=32'h000C007A;
14'd7251:data <=32'h0022007A;14'd7252:data <=32'h00370073;14'd7253:data <=32'h00470067;
14'd7254:data <=32'h00520055;14'd7255:data <=32'h00560045;14'd7256:data <=32'h00560037;
14'd7257:data <=32'h0056002B;14'd7258:data <=32'h00540024;14'd7259:data <=32'h0053001C;
14'd7260:data <=32'h00540015;14'd7261:data <=32'h0052000C;14'd7262:data <=32'h00510003;
14'd7263:data <=32'h004DFFFC;14'd7264:data <=32'h0046FFF4;14'd7265:data <=32'h003FFFF0;
14'd7266:data <=32'h0038FFED;14'd7267:data <=32'h0033FFEC;14'd7268:data <=32'h002EFFEB;
14'd7269:data <=32'h002AFFEB;14'd7270:data <=32'h0026FFEB;14'd7271:data <=32'h001FFFEB;
14'd7272:data <=32'h0018FFEE;14'd7273:data <=32'h0011FFF6;14'd7274:data <=32'h000D0003;
14'd7275:data <=32'h000F0013;14'd7276:data <=32'h001A0024;14'd7277:data <=32'h002D0031;
14'd7278:data <=32'h004A0037;14'd7279:data <=32'h006A0033;14'd7280:data <=32'h00890021;
14'd7281:data <=32'h00A40005;14'd7282:data <=32'h00B7FFE0;14'd7283:data <=32'h00BDFFB4;
14'd7284:data <=32'h00B7FF87;14'd7285:data <=32'h00A7FF5C;14'd7286:data <=32'h008DFF34;
14'd7287:data <=32'h0069FF10;14'd7288:data <=32'h003CFEF7;14'd7289:data <=32'h0009FEE6;
14'd7290:data <=32'hFFD0FEE0;14'd7291:data <=32'hFF97FEEA;14'd7292:data <=32'hFF60FF02;
14'd7293:data <=32'hFF30FF29;14'd7294:data <=32'hFF0EFF5B;14'd7295:data <=32'hFEFDFF92;
14'd7296:data <=32'hFF58FF8E;14'd7297:data <=32'hFF3CFFA2;14'd7298:data <=32'hFF22FFAE;
14'd7299:data <=32'hFF0AFF9F;14'd7300:data <=32'hFF40FFD4;14'd7301:data <=32'hFF40FFE9;
14'd7302:data <=32'hFF40FFFC;14'd7303:data <=32'hFF400012;14'd7304:data <=32'hFF45002B;
14'd7305:data <=32'hFF4E0043;14'd7306:data <=32'hFF5B005A;14'd7307:data <=32'hFF6D006D;
14'd7308:data <=32'hFF7F007C;14'd7309:data <=32'hFF930088;14'd7310:data <=32'hFFA80092;
14'd7311:data <=32'hFFBD009A;14'd7312:data <=32'hFFD6009F;14'd7313:data <=32'hFFF100A0;
14'd7314:data <=32'h000D009B;14'd7315:data <=32'h0028008E;14'd7316:data <=32'h003E0077;
14'd7317:data <=32'h004A005D;14'd7318:data <=32'h004D0040;14'd7319:data <=32'h00470027;
14'd7320:data <=32'h00370014;14'd7321:data <=32'h0026000B;14'd7322:data <=32'h00140009;
14'd7323:data <=32'h00050010;14'd7324:data <=32'hFFFD001B;14'd7325:data <=32'hFFFA0026;
14'd7326:data <=32'hFFFD0031;14'd7327:data <=32'h0001003A;14'd7328:data <=32'h000A0041;
14'd7329:data <=32'h00140045;14'd7330:data <=32'h001F0047;14'd7331:data <=32'h002B0046;
14'd7332:data <=32'h00380042;14'd7333:data <=32'h00420039;14'd7334:data <=32'h004A002D;
14'd7335:data <=32'h004D001E;14'd7336:data <=32'h00480011;14'd7337:data <=32'h00400007;
14'd7338:data <=32'h00350003;14'd7339:data <=32'h002A0007;14'd7340:data <=32'h00220010;
14'd7341:data <=32'h0022001F;14'd7342:data <=32'h002B002D;14'd7343:data <=32'h003C0037;
14'd7344:data <=32'h0052003A;14'd7345:data <=32'h00690035;14'd7346:data <=32'h007F0027;
14'd7347:data <=32'h00900013;14'd7348:data <=32'h009CFFFB;14'd7349:data <=32'h00A4FFE0;
14'd7350:data <=32'h00A4FFC5;14'd7351:data <=32'h00A0FFA9;14'd7352:data <=32'h0098FF8C;
14'd7353:data <=32'h0089FF71;14'd7354:data <=32'h0074FF58;14'd7355:data <=32'h0059FF42;
14'd7356:data <=32'h0039FF35;14'd7357:data <=32'h0017FF2F;14'd7358:data <=32'hFFF7FF33;
14'd7359:data <=32'hFFDBFF3B;14'd7360:data <=32'hFFBAFEFB;14'd7361:data <=32'hFF87FF01;
14'd7362:data <=32'hFF70FF15;14'd7363:data <=32'hFFD9FF31;14'd7364:data <=32'hFFF9FF40;
14'd7365:data <=32'hFFDBFF32;14'd7366:data <=32'hFFB6FF2C;14'd7367:data <=32'hFF8CFF2E;
14'd7368:data <=32'hFF61FF3E;14'd7369:data <=32'hFF3AFF5B;14'd7370:data <=32'hFF1CFF80;
14'd7371:data <=32'hFF08FFAC;14'd7372:data <=32'hFEFCFFDB;14'd7373:data <=32'hFEFC000A;
14'd7374:data <=32'hFF040039;14'd7375:data <=32'hFF170066;14'd7376:data <=32'hFF35008E;
14'd7377:data <=32'hFF5C00AF;14'd7378:data <=32'hFF8A00C5;14'd7379:data <=32'hFFBC00CD;
14'd7380:data <=32'hFFEF00C5;14'd7381:data <=32'h001A00B0;14'd7382:data <=32'h003A008F;
14'd7383:data <=32'h004C006A;14'd7384:data <=32'h004F0044;14'd7385:data <=32'h00480024;
14'd7386:data <=32'h0039000C;14'd7387:data <=32'h0025FFFD;14'd7388:data <=32'h0012FFF6;
14'd7389:data <=32'h0000FFF5;14'd7390:data <=32'hFFEFFFF8;14'd7391:data <=32'hFFE2FFFF;
14'd7392:data <=32'hFFD7000A;14'd7393:data <=32'hFFCF0016;14'd7394:data <=32'hFFCA0024;
14'd7395:data <=32'hFFCA0036;14'd7396:data <=32'hFFD00046;14'd7397:data <=32'hFFD90054;
14'd7398:data <=32'hFFE7005E;14'd7399:data <=32'hFFF60064;14'd7400:data <=32'h00040066;
14'd7401:data <=32'h000F0065;14'd7402:data <=32'h00190065;14'd7403:data <=32'h00210065;
14'd7404:data <=32'h002A0068;14'd7405:data <=32'h0037006A;14'd7406:data <=32'h0048006B;
14'd7407:data <=32'h005C0069;14'd7408:data <=32'h0071005F;14'd7409:data <=32'h0084004F;
14'd7410:data <=32'h00940039;14'd7411:data <=32'h009C001F;14'd7412:data <=32'h009D0004;
14'd7413:data <=32'h0096FFEC;14'd7414:data <=32'h008CFFD9;14'd7415:data <=32'h007EFFCC;
14'd7416:data <=32'h0072FFC2;14'd7417:data <=32'h0067FFBD;14'd7418:data <=32'h005CFFB8;
14'd7419:data <=32'h0053FFB5;14'd7420:data <=32'h004BFFB5;14'd7421:data <=32'h0045FFB5;
14'd7422:data <=32'h0043FFB8;14'd7423:data <=32'h0046FFB9;14'd7424:data <=32'h0089FF3C;
14'd7425:data <=32'h006CFF1E;14'd7426:data <=32'h0046FF1D;14'd7427:data <=32'h004EFF9D;
14'd7428:data <=32'h0089FFA0;14'd7429:data <=32'h0086FF79;14'd7430:data <=32'h0076FF52;
14'd7431:data <=32'h0058FF2D;14'd7432:data <=32'h002EFF14;14'd7433:data <=32'hFFFEFF08;
14'd7434:data <=32'hFFCDFF08;14'd7435:data <=32'hFF9EFF13;14'd7436:data <=32'hFF74FF29;
14'd7437:data <=32'hFF50FF47;14'd7438:data <=32'hFF32FF6B;14'd7439:data <=32'hFF1CFF96;
14'd7440:data <=32'hFF11FFC6;14'd7441:data <=32'hFF11FFF7;14'd7442:data <=32'hFF1F0026;
14'd7443:data <=32'hFF39004E;14'd7444:data <=32'hFF5B006C;14'd7445:data <=32'hFF82007D;
14'd7446:data <=32'hFFA80082;14'd7447:data <=32'hFFC9007C;14'd7448:data <=32'hFFE20070;
14'd7449:data <=32'hFFF40061;14'd7450:data <=32'h00010052;14'd7451:data <=32'h00080044;
14'd7452:data <=32'h000E0037;14'd7453:data <=32'h0012002A;14'd7454:data <=32'h0013001E;
14'd7455:data <=32'h0013000F;14'd7456:data <=32'h000D0000;14'd7457:data <=32'h0003FFF3;
14'd7458:data <=32'hFFF4FFEA;14'd7459:data <=32'hFFE2FFE7;14'd7460:data <=32'hFFCFFFE8;
14'd7461:data <=32'hFFBEFFF0;14'd7462:data <=32'hFFAEFFFD;14'd7463:data <=32'hFFA3000D;
14'd7464:data <=32'hFF9A0020;14'd7465:data <=32'hFF940036;14'd7466:data <=32'hFF92004E;
14'd7467:data <=32'hFF960069;14'd7468:data <=32'hFFA00087;14'd7469:data <=32'hFFB300A4;
14'd7470:data <=32'hFFD100BC;14'd7471:data <=32'hFFF600CF;14'd7472:data <=32'h002300D6;
14'd7473:data <=32'h005000D1;14'd7474:data <=32'h007A00BD;14'd7475:data <=32'h009C009E;
14'd7476:data <=32'h00B40078;14'd7477:data <=32'h00BF0050;14'd7478:data <=32'h00BE002A;
14'd7479:data <=32'h00B40009;14'd7480:data <=32'h00A6FFEF;14'd7481:data <=32'h0095FFDB;
14'd7482:data <=32'h0081FFCF;14'd7483:data <=32'h006CFFC7;14'd7484:data <=32'h005CFFC5;
14'd7485:data <=32'h004CFFCA;14'd7486:data <=32'h0041FFD3;14'd7487:data <=32'h003EFFDF;
14'd7488:data <=32'h0080FFEF;14'd7489:data <=32'h008FFFE2;14'd7490:data <=32'h0089FFCA;
14'd7491:data <=32'h004DFFC0;14'd7492:data <=32'h0088FFD3;14'd7493:data <=32'h008EFFBB;
14'd7494:data <=32'h008CFF9E;14'd7495:data <=32'h0080FF82;14'd7496:data <=32'h006BFF6A;
14'd7497:data <=32'h0050FF59;14'd7498:data <=32'h0034FF50;14'd7499:data <=32'h0017FF4F;
14'd7500:data <=32'hFFFEFF51;14'd7501:data <=32'hFFE7FF57;14'd7502:data <=32'hFFD1FF5F;
14'd7503:data <=32'hFFBDFF6A;14'd7504:data <=32'hFFAAFF79;14'd7505:data <=32'hFF9AFF8B;
14'd7506:data <=32'hFF90FFA0;14'd7507:data <=32'hFF8CFFB5;14'd7508:data <=32'hFF8CFFCA;
14'd7509:data <=32'hFF92FFD9;14'd7510:data <=32'hFF98FFE3;14'd7511:data <=32'hFF9BFFEB;
14'd7512:data <=32'hFF9CFFF1;14'd7513:data <=32'hFF9BFFF9;14'd7514:data <=32'hFF9A0004;
14'd7515:data <=32'hFF9B0012;14'd7516:data <=32'hFFA20022;14'd7517:data <=32'hFFAE0032;
14'd7518:data <=32'hFFC0003D;14'd7519:data <=32'hFFD50040;14'd7520:data <=32'hFFEB003C;
14'd7521:data <=32'hFFFD0030;14'd7522:data <=32'h0008001F;14'd7523:data <=32'h000D000C;
14'd7524:data <=32'h000BFFF8;14'd7525:data <=32'h0002FFE6;14'd7526:data <=32'hFFF4FFD6;
14'd7527:data <=32'hFFE1FFCC;14'd7528:data <=32'hFFCBFFC7;14'd7529:data <=32'hFFB1FFC8;
14'd7530:data <=32'hFF96FFD1;14'd7531:data <=32'hFF7BFFE3;14'd7532:data <=32'hFF65FFFE;
14'd7533:data <=32'hFF550022;14'd7534:data <=32'hFF52004C;14'd7535:data <=32'hFF5C0077;
14'd7536:data <=32'hFF71009F;14'd7537:data <=32'hFF9300BE;14'd7538:data <=32'hFFBB00D1;
14'd7539:data <=32'hFFE500DA;14'd7540:data <=32'h000C00D7;14'd7541:data <=32'h002F00CA;
14'd7542:data <=32'h004A00BB;14'd7543:data <=32'h006000A9;14'd7544:data <=32'h00710095;
14'd7545:data <=32'h007E0083;14'd7546:data <=32'h008A0071;14'd7547:data <=32'h0092005D;
14'd7548:data <=32'h0097004A;14'd7549:data <=32'h00990038;14'd7550:data <=32'h00990027;
14'd7551:data <=32'h0097001A;14'd7552:data <=32'h0030FFFD;14'd7553:data <=32'h00350012;
14'd7554:data <=32'h004E001A;14'd7555:data <=32'h00B2FFF1;14'd7556:data <=32'h00E6FFF2;
14'd7557:data <=32'h00E3FFC9;14'd7558:data <=32'h00D4FFA1;14'd7559:data <=32'h00BBFF7B;
14'd7560:data <=32'h0097FF5F;14'd7561:data <=32'h006EFF51;14'd7562:data <=32'h0046FF4E;
14'd7563:data <=32'h0021FF56;14'd7564:data <=32'h0006FF66;14'd7565:data <=32'hFFF2FF7A;
14'd7566:data <=32'hFFE6FF8E;14'd7567:data <=32'hFFE1FFA1;14'd7568:data <=32'hFFE0FFB1;
14'd7569:data <=32'hFFE2FFBF;14'd7570:data <=32'hFFE8FFC9;14'd7571:data <=32'hFFF0FFD0;
14'd7572:data <=32'hFFF9FFD2;14'd7573:data <=32'h0002FFCE;14'd7574:data <=32'h0009FFC4;
14'd7575:data <=32'h0009FFB6;14'd7576:data <=32'h0001FFA7;14'd7577:data <=32'hFFF2FF9C;
14'd7578:data <=32'hFFDDFF97;14'd7579:data <=32'hFFC5FF9C;14'd7580:data <=32'hFFB0FFA9;
14'd7581:data <=32'hFFA1FFBD;14'd7582:data <=32'hFF9BFFD4;14'd7583:data <=32'hFF9DFFEA;
14'd7584:data <=32'hFFA7FFFD;14'd7585:data <=32'hFFB50009;14'd7586:data <=32'hFFC4000F;
14'd7587:data <=32'hFFD10010;14'd7588:data <=32'hFFDD000D;14'd7589:data <=32'hFFE60007;
14'd7590:data <=32'hFFEDFFFF;14'd7591:data <=32'hFFF0FFF4;14'd7592:data <=32'hFFEFFFE7;
14'd7593:data <=32'hFFE9FFDA;14'd7594:data <=32'hFFDEFFCF;14'd7595:data <=32'hFFCEFFC8;
14'd7596:data <=32'hFFBAFFC5;14'd7597:data <=32'hFFA4FFCA;14'd7598:data <=32'hFF90FFD7;
14'd7599:data <=32'hFF80FFE9;14'd7600:data <=32'hFF77FFFF;14'd7601:data <=32'hFF720017;
14'd7602:data <=32'hFF75002C;14'd7603:data <=32'hFF7A003E;14'd7604:data <=32'hFF80004D;
14'd7605:data <=32'hFF85005B;14'd7606:data <=32'hFF87006A;14'd7607:data <=32'hFF8C007D;
14'd7608:data <=32'hFF940094;14'd7609:data <=32'hFFA100AC;14'd7610:data <=32'hFFB600C5;
14'd7611:data <=32'hFFD200D9;14'd7612:data <=32'hFFF500E9;14'd7613:data <=32'h001B00F0;
14'd7614:data <=32'h004300EF;14'd7615:data <=32'h006C00E8;14'd7616:data <=32'h004B0020;
14'd7617:data <=32'h0042002E;14'd7618:data <=32'h0044004F;14'd7619:data <=32'h00A200C7;
14'd7620:data <=32'h00FC00C3;14'd7621:data <=32'h011F008C;14'd7622:data <=32'h012F004B;
14'd7623:data <=32'h0130000A;14'd7624:data <=32'h011DFFCB;14'd7625:data <=32'h00FAFF97;
14'd7626:data <=32'h00CEFF72;14'd7627:data <=32'h009EFF5D;14'd7628:data <=32'h006FFF57;
14'd7629:data <=32'h0047FF5C;14'd7630:data <=32'h0026FF69;14'd7631:data <=32'h000CFF7A;
14'd7632:data <=32'hFFF9FF8F;14'd7633:data <=32'hFFEDFFA3;14'd7634:data <=32'hFFE7FFBA;
14'd7635:data <=32'hFFE9FFCE;14'd7636:data <=32'hFFF2FFE0;14'd7637:data <=32'h0000FFEA;
14'd7638:data <=32'h0010FFED;14'd7639:data <=32'h001EFFEA;14'd7640:data <=32'h0028FFDE;
14'd7641:data <=32'h002BFFCF;14'd7642:data <=32'h0027FFC0;14'd7643:data <=32'h001DFFB4;
14'd7644:data <=32'h0011FFAE;14'd7645:data <=32'h0004FFAD;14'd7646:data <=32'hFFF9FFB1;
14'd7647:data <=32'hFFF3FFB6;14'd7648:data <=32'hFFEFFFBB;14'd7649:data <=32'hFFEDFFBD;
14'd7650:data <=32'hFFECFFBE;14'd7651:data <=32'hFFE8FFBC;14'd7652:data <=32'hFFE2FFBA;
14'd7653:data <=32'hFFDAFFBB;14'd7654:data <=32'hFFD3FFBF;14'd7655:data <=32'hFFCBFFC4;
14'd7656:data <=32'hFFC8FFCB;14'd7657:data <=32'hFFC4FFD1;14'd7658:data <=32'hFFC3FFD6;
14'd7659:data <=32'hFFC1FFDB;14'd7660:data <=32'hFFC0FFDE;14'd7661:data <=32'hFFBFFFE2;
14'd7662:data <=32'hFFBEFFE6;14'd7663:data <=32'hFFBEFFEA;14'd7664:data <=32'hFFC1FFEE;
14'd7665:data <=32'hFFC4FFEE;14'd7666:data <=32'hFFC7FFEB;14'd7667:data <=32'hFFC7FFE3;
14'd7668:data <=32'hFFC0FFD8;14'd7669:data <=32'hFFB1FFCD;14'd7670:data <=32'hFF9AFFC8;
14'd7671:data <=32'hFF7CFFCC;14'd7672:data <=32'hFF5DFFDC;14'd7673:data <=32'hFF41FFF7;
14'd7674:data <=32'hFF2C001F;14'd7675:data <=32'hFF23004E;14'd7676:data <=32'hFF270080;
14'd7677:data <=32'hFF3800B0;14'd7678:data <=32'hFF5400DC;14'd7679:data <=32'hFF7B0103;
14'd7680:data <=32'hFFDE008B;14'd7681:data <=32'hFFE400A4;14'd7682:data <=32'hFFDC00BA;
14'd7683:data <=32'hFFB50101;14'd7684:data <=32'h001C012E;14'd7685:data <=32'h00570120;
14'd7686:data <=32'h008B0103;14'd7687:data <=32'h00B500DA;14'd7688:data <=32'h00D200AA;
14'd7689:data <=32'h00DE0079;14'd7690:data <=32'h00DE004B;14'd7691:data <=32'h00D50024;
14'd7692:data <=32'h00C60005;14'd7693:data <=32'h00B6FFED;14'd7694:data <=32'h00A6FFDA;
14'd7695:data <=32'h0096FFCB;14'd7696:data <=32'h0085FFBC;14'd7697:data <=32'h0072FFB3;
14'd7698:data <=32'h005FFFAB;14'd7699:data <=32'h004BFFA8;14'd7700:data <=32'h003AFFAA;
14'd7701:data <=32'h002DFFB0;14'd7702:data <=32'h0023FFB6;14'd7703:data <=32'h001CFFBC;
14'd7704:data <=32'h0017FFC1;14'd7705:data <=32'h0010FFC4;14'd7706:data <=32'h000AFFC7;
14'd7707:data <=32'h0003FFCE;14'd7708:data <=32'hFFFFFFD7;14'd7709:data <=32'hFFFDFFE3;
14'd7710:data <=32'h0002FFF0;14'd7711:data <=32'h000DFFFA;14'd7712:data <=32'h001CFFFE;
14'd7713:data <=32'h002EFFFB;14'd7714:data <=32'h003CFFF0;14'd7715:data <=32'h0047FFDD;
14'd7716:data <=32'h004AFFC7;14'd7717:data <=32'h0044FFB1;14'd7718:data <=32'h0037FF9F;
14'd7719:data <=32'h0027FF91;14'd7720:data <=32'h0013FF88;14'd7721:data <=32'hFFFFFF84;
14'd7722:data <=32'hFFEBFF87;14'd7723:data <=32'hFFD9FF8C;14'd7724:data <=32'hFFC9FF96;
14'd7725:data <=32'hFFBBFFA3;14'd7726:data <=32'hFFB2FFB2;14'd7727:data <=32'hFFAEFFC3;
14'd7728:data <=32'hFFB0FFD3;14'd7729:data <=32'hFFB7FFE0;14'd7730:data <=32'hFFC3FFE7;
14'd7731:data <=32'hFFD0FFE5;14'd7732:data <=32'hFFDAFFDC;14'd7733:data <=32'hFFDDFFCC;
14'd7734:data <=32'hFFD5FFBA;14'd7735:data <=32'hFFC4FFA9;14'd7736:data <=32'hFFAAFFA1;
14'd7737:data <=32'hFF89FFA2;14'd7738:data <=32'hFF69FFAF;14'd7739:data <=32'hFF4DFFC7;
14'd7740:data <=32'hFF38FFE6;14'd7741:data <=32'hFF2C000A;14'd7742:data <=32'hFF280031;
14'd7743:data <=32'hFF2A0058;14'd7744:data <=32'hFF2D001C;14'd7745:data <=32'hFF160051;
14'd7746:data <=32'hFF150077;14'd7747:data <=32'hFF4F0065;14'd7748:data <=32'hFF9100A3;
14'd7749:data <=32'hFFAD00AF;14'd7750:data <=32'hFFC900B2;14'd7751:data <=32'hFFE400B1;
14'd7752:data <=32'hFFFA00A9;14'd7753:data <=32'h000900A0;14'd7754:data <=32'h00140099;
14'd7755:data <=32'h001D0095;14'd7756:data <=32'h00270097;14'd7757:data <=32'h00360098;
14'd7758:data <=32'h004B0098;14'd7759:data <=32'h00630092;14'd7760:data <=32'h007C0085;
14'd7761:data <=32'h00910070;14'd7762:data <=32'h00A20055;14'd7763:data <=32'h00AB0037;
14'd7764:data <=32'h00AD0019;14'd7765:data <=32'h00A9FFFB;14'd7766:data <=32'h009FFFE0;
14'd7767:data <=32'h0091FFC7;14'd7768:data <=32'h007DFFB2;14'd7769:data <=32'h0065FFA1;
14'd7770:data <=32'h0048FF97;14'd7771:data <=32'h0029FF96;14'd7772:data <=32'h000AFF9E;
14'd7773:data <=32'hFFF1FFB1;14'd7774:data <=32'hFFE0FFCB;14'd7775:data <=32'hFFDBFFEA;
14'd7776:data <=32'hFFE10007;14'd7777:data <=32'hFFF2001D;14'd7778:data <=32'h000A002B;
14'd7779:data <=32'h0025002F;14'd7780:data <=32'h003D0029;14'd7781:data <=32'h0051001B;
14'd7782:data <=32'h00600009;14'd7783:data <=32'h006AFFF4;14'd7784:data <=32'h006CFFE0;
14'd7785:data <=32'h006BFFCC;14'd7786:data <=32'h0066FFB8;14'd7787:data <=32'h005DFFA5;
14'd7788:data <=32'h0051FF95;14'd7789:data <=32'h0041FF87;14'd7790:data <=32'h002EFF7D;
14'd7791:data <=32'h001BFF78;14'd7792:data <=32'h0009FF78;14'd7793:data <=32'hFFF9FF7B;
14'd7794:data <=32'hFFEDFF7F;14'd7795:data <=32'hFFE5FF82;14'd7796:data <=32'hFFDCFF82;
14'd7797:data <=32'hFFD3FF7F;14'd7798:data <=32'hFFC5FF7B;14'd7799:data <=32'hFFB1FF78;
14'd7800:data <=32'hFF9AFF7B;14'd7801:data <=32'hFF81FF85;14'd7802:data <=32'hFF68FF97;
14'd7803:data <=32'hFF56FFB1;14'd7804:data <=32'hFF49FFCE;14'd7805:data <=32'hFF47FFED;
14'd7806:data <=32'hFF4A0009;14'd7807:data <=32'hFF540021;14'd7808:data <=32'hFF6AFF63;
14'd7809:data <=32'hFF28FF79;14'd7810:data <=32'hFF04FFAD;14'd7811:data <=32'hFF6B002B;
14'd7812:data <=32'hFFA7005B;14'd7813:data <=32'hFFB90057;14'd7814:data <=32'hFFC9004E;
14'd7815:data <=32'hFFD10043;14'd7816:data <=32'hFFD30035;14'd7817:data <=32'hFFCA002B;
14'd7818:data <=32'hFFBC0028;14'd7819:data <=32'hFFAC002F;14'd7820:data <=32'hFF9D0040;
14'd7821:data <=32'hFF98005B;14'd7822:data <=32'hFF9C007A;14'd7823:data <=32'hFFAD0097;
14'd7824:data <=32'hFFC800AF;14'd7825:data <=32'hFFEB00BE;14'd7826:data <=32'h001000C1;
14'd7827:data <=32'h003300BC;14'd7828:data <=32'h005500AE;14'd7829:data <=32'h00720099;
14'd7830:data <=32'h0089007F;14'd7831:data <=32'h009B0061;14'd7832:data <=32'h00A40040;
14'd7833:data <=32'h00A5001B;14'd7834:data <=32'h009CFFF9;14'd7835:data <=32'h0089FFDA;
14'd7836:data <=32'h006FFFC3;14'd7837:data <=32'h0050FFB6;14'd7838:data <=32'h0031FFB6;
14'd7839:data <=32'h0016FFBF;14'd7840:data <=32'h0003FFD0;14'd7841:data <=32'hFFF8FFE4;
14'd7842:data <=32'hFFF5FFF8;14'd7843:data <=32'hFFF80008;14'd7844:data <=32'hFFFF0015;
14'd7845:data <=32'h0007001F;14'd7846:data <=32'h00110026;14'd7847:data <=32'h001B002D;
14'd7848:data <=32'h00260032;14'd7849:data <=32'h00350036;14'd7850:data <=32'h00460037;
14'd7851:data <=32'h005A0033;14'd7852:data <=32'h0070002A;14'd7853:data <=32'h0083001B;
14'd7854:data <=32'h00920005;14'd7855:data <=32'h009EFFEC;14'd7856:data <=32'h00A3FFD1;
14'd7857:data <=32'h00A5FFB3;14'd7858:data <=32'h00A0FF95;14'd7859:data <=32'h0096FF75;
14'd7860:data <=32'h0087FF55;14'd7861:data <=32'h0070FF36;14'd7862:data <=32'h0050FF1A;
14'd7863:data <=32'h0025FF02;14'd7864:data <=32'hFFF3FEF5;14'd7865:data <=32'hFFBCFEF8;
14'd7866:data <=32'hFF87FF08;14'd7867:data <=32'hFF59FF28;14'd7868:data <=32'hFF35FF54;
14'd7869:data <=32'hFF20FF84;14'd7870:data <=32'hFF19FFB5;14'd7871:data <=32'hFF20FFE2;
14'd7872:data <=32'hFFD9FF69;14'd7873:data <=32'hFFABFF58;14'd7874:data <=32'hFF6DFF63;
14'd7875:data <=32'hFF2AFFEC;14'd7876:data <=32'hFF670030;14'd7877:data <=32'hFF81003C;
14'd7878:data <=32'hFF9B0040;14'd7879:data <=32'hFFB1003B;14'd7880:data <=32'hFFC00030;
14'd7881:data <=32'hFFC60021;14'd7882:data <=32'hFFC30013;14'd7883:data <=32'hFFB7000B;
14'd7884:data <=32'hFFA8000C;14'd7885:data <=32'hFF990017;14'd7886:data <=32'hFF8F0029;
14'd7887:data <=32'hFF8D0040;14'd7888:data <=32'hFF940058;14'd7889:data <=32'hFFA2006C;
14'd7890:data <=32'hFFB50079;14'd7891:data <=32'hFFC90082;14'd7892:data <=32'hFFDC0087;
14'd7893:data <=32'hFFF00088;14'd7894:data <=32'h00020087;14'd7895:data <=32'h00160082;
14'd7896:data <=32'h0027007B;14'd7897:data <=32'h0038006E;14'd7898:data <=32'h0045005E;
14'd7899:data <=32'h004D004C;14'd7900:data <=32'h0050003B;14'd7901:data <=32'h004B002A;
14'd7902:data <=32'h0046001E;14'd7903:data <=32'h003D0017;14'd7904:data <=32'h00370013;
14'd7905:data <=32'h00340010;14'd7906:data <=32'h0031000D;14'd7907:data <=32'h002F0009;
14'd7908:data <=32'h002B0003;14'd7909:data <=32'h0023FFFD;14'd7910:data <=32'h0018FFFA;
14'd7911:data <=32'h000BFFFC;14'd7912:data <=32'hFFFE0006;14'd7913:data <=32'hFFF30015;
14'd7914:data <=32'hFFF00029;14'd7915:data <=32'hFFF50040;14'd7916:data <=32'h00030057;
14'd7917:data <=32'h00190068;14'd7918:data <=32'h00360073;14'd7919:data <=32'h00560076;
14'd7920:data <=32'h00780071;14'd7921:data <=32'h009B0063;14'd7922:data <=32'h00BB004C;
14'd7923:data <=32'h00D8002C;14'd7924:data <=32'h00EE0004;14'd7925:data <=32'h00FCFFD2;
14'd7926:data <=32'h00FCFF9B;14'd7927:data <=32'h00EDFF63;14'd7928:data <=32'h00CDFF2D;
14'd7929:data <=32'h00A0FF02;14'd7930:data <=32'h0067FEE5;14'd7931:data <=32'h002BFED9;
14'd7932:data <=32'hFFEFFEDF;14'd7933:data <=32'hFFBBFEF2;14'd7934:data <=32'hFF90FF10;
14'd7935:data <=32'hFF72FF32;14'd7936:data <=32'hFFD4FF5C;14'd7937:data <=32'hFFB9FF52;
14'd7938:data <=32'hFF97FF42;14'd7939:data <=32'hFF69FF2A;14'd7940:data <=32'hFF7DFF70;
14'd7941:data <=32'hFF72FF86;14'd7942:data <=32'hFF6CFF9B;14'd7943:data <=32'hFF68FFB1;
14'd7944:data <=32'hFF67FFC2;14'd7945:data <=32'hFF67FFD1;14'd7946:data <=32'hFF65FFDE;
14'd7947:data <=32'hFF60FFED;14'd7948:data <=32'hFF5D0000;14'd7949:data <=32'hFF5B0017;
14'd7950:data <=32'hFF600030;14'd7951:data <=32'hFF6D004A;14'd7952:data <=32'hFF820060;
14'd7953:data <=32'hFF9C006F;14'd7954:data <=32'hFFB90074;14'd7955:data <=32'hFFD20070;
14'd7956:data <=32'hFFE60065;14'd7957:data <=32'hFFF40057;14'd7958:data <=32'hFFFB004A;
14'd7959:data <=32'hFFFE003E;14'd7960:data <=32'hFFFD0035;14'd7961:data <=32'hFFFC002E;
14'd7962:data <=32'hFFF80029;14'd7963:data <=32'hFFF30026;14'd7964:data <=32'hFFED0025;
14'd7965:data <=32'hFFE60028;14'd7966:data <=32'hFFE2002F;14'd7967:data <=32'hFFE10039;
14'd7968:data <=32'hFFE40045;14'd7969:data <=32'hFFEE0050;14'd7970:data <=32'hFFFC0056;
14'd7971:data <=32'h000C0057;14'd7972:data <=32'h001D0051;14'd7973:data <=32'h00280044;
14'd7974:data <=32'h002D0034;14'd7975:data <=32'h002A0024;14'd7976:data <=32'h00210018;
14'd7977:data <=32'h00120014;14'd7978:data <=32'h00040018;14'd7979:data <=32'hFFFA0022;
14'd7980:data <=32'hFFF3002F;14'd7981:data <=32'hFFF30041;14'd7982:data <=32'hFFFA0053;
14'd7983:data <=32'h00070064;14'd7984:data <=32'h00180071;14'd7985:data <=32'h002E007B;
14'd7986:data <=32'h00480081;14'd7987:data <=32'h00660080;14'd7988:data <=32'h00840077;
14'd7989:data <=32'h00A40065;14'd7990:data <=32'h00C1004A;14'd7991:data <=32'h00D50027;
14'd7992:data <=32'h00E0FFFD;14'd7993:data <=32'h00DEFFD4;14'd7994:data <=32'h00D2FFAC;
14'd7995:data <=32'h00BDFF8B;14'd7996:data <=32'h00A4FF73;14'd7997:data <=32'h008BFF63;
14'd7998:data <=32'h0074FF58;14'd7999:data <=32'h0060FF4E;14'd8000:data <=32'h004AFF18;
14'd8001:data <=32'h0025FF04;14'd8002:data <=32'h000FFEFF;14'd8003:data <=32'h0061FF25;
14'd8004:data <=32'h006DFF3D;14'd8005:data <=32'h0051FF27;14'd8006:data <=32'h002EFF15;
14'd8007:data <=32'h0007FF0A;14'd8008:data <=32'hFFDFFF08;14'd8009:data <=32'hFFB6FF0C;
14'd8010:data <=32'hFF8BFF17;14'd8011:data <=32'hFF62FF2D;14'd8012:data <=32'hFF3CFF4C;
14'd8013:data <=32'hFF1CFF78;14'd8014:data <=32'hFF09FFAB;14'd8015:data <=32'hFF04FFE3;
14'd8016:data <=32'hFF100019;14'd8017:data <=32'hFF2C0048;14'd8018:data <=32'hFF510069;
14'd8019:data <=32'hFF7B007E;14'd8020:data <=32'hFFA60083;14'd8021:data <=32'hFFCB007D;
14'd8022:data <=32'hFFE9006F;14'd8023:data <=32'hFFFF005C;14'd8024:data <=32'h000E0047;
14'd8025:data <=32'h00150031;14'd8026:data <=32'h0016001B;14'd8027:data <=32'h00110008;
14'd8028:data <=32'h0007FFF7;14'd8029:data <=32'hFFF6FFEC;14'd8030:data <=32'hFFE3FFE6;
14'd8031:data <=32'hFFCEFFEA;14'd8032:data <=32'hFFBEFFF4;14'd8033:data <=32'hFFB30004;
14'd8034:data <=32'hFFAF0017;14'd8035:data <=32'hFFB20029;14'd8036:data <=32'hFFB90036;
14'd8037:data <=32'hFFC3003E;14'd8038:data <=32'hFFCD0043;14'd8039:data <=32'hFFD30045;
14'd8040:data <=32'hFFD50047;14'd8041:data <=32'hFFD7004A;14'd8042:data <=32'hFFD80050;
14'd8043:data <=32'hFFDC005A;14'd8044:data <=32'hFFE20065;14'd8045:data <=32'hFFED006E;
14'd8046:data <=32'hFFFC0076;14'd8047:data <=32'h000C007A;14'd8048:data <=32'h001D007A;
14'd8049:data <=32'h002D0076;14'd8050:data <=32'h003A0071;14'd8051:data <=32'h0047006B;
14'd8052:data <=32'h00530063;14'd8053:data <=32'h005E005A;14'd8054:data <=32'h0069004F;
14'd8055:data <=32'h00710040;14'd8056:data <=32'h00760031;14'd8057:data <=32'h00760023;
14'd8058:data <=32'h00720018;14'd8059:data <=32'h006C0011;14'd8060:data <=32'h00690010;
14'd8061:data <=32'h006A0014;14'd8062:data <=32'h00740017;14'd8063:data <=32'h00840015;
14'd8064:data <=32'h00DDFFAA;14'd8065:data <=32'h00D9FF80;14'd8066:data <=32'h00C0FF6F;
14'd8067:data <=32'h00A6FFE4;14'd8068:data <=32'h00D9FFF4;14'd8069:data <=32'h00E1FFC8;
14'd8070:data <=32'h00DFFF9B;14'd8071:data <=32'h00D0FF6F;14'd8072:data <=32'h00B9FF44;
14'd8073:data <=32'h0098FF1F;14'd8074:data <=32'h006EFF01;14'd8075:data <=32'h003AFEEB;
14'd8076:data <=32'h0002FEE2;14'd8077:data <=32'hFFC7FEEA;14'd8078:data <=32'hFF90FF02;
14'd8079:data <=32'hFF62FF28;14'd8080:data <=32'hFF42FF58;14'd8081:data <=32'hFF33FF8B;
14'd8082:data <=32'hFF33FFBD;14'd8083:data <=32'hFF3EFFE7;14'd8084:data <=32'hFF530009;
14'd8085:data <=32'hFF6A0022;14'd8086:data <=32'hFF820033;14'd8087:data <=32'hFF9A003C;
14'd8088:data <=32'hFFB10042;14'd8089:data <=32'hFFC60043;14'd8090:data <=32'hFFDB0040;
14'd8091:data <=32'hFFEE0037;14'd8092:data <=32'hFFFD002A;14'd8093:data <=32'h0006001A;
14'd8094:data <=32'h00090008;14'd8095:data <=32'h0006FFF7;14'd8096:data <=32'hFFFEFFEA;
14'd8097:data <=32'hFFF4FFE2;14'd8098:data <=32'hFFE9FFDC;14'd8099:data <=32'hFFDEFFD9;
14'd8100:data <=32'hFFD3FFD6;14'd8101:data <=32'hFFC7FFD5;14'd8102:data <=32'hFFB9FFD5;
14'd8103:data <=32'hFFA8FFD8;14'd8104:data <=32'hFF95FFE1;14'd8105:data <=32'hFF81FFF0;
14'd8106:data <=32'hFF700008;14'd8107:data <=32'hFF650026;14'd8108:data <=32'hFF640049;
14'd8109:data <=32'hFF6E006C;14'd8110:data <=32'hFF81008D;14'd8111:data <=32'hFF9E00A6;
14'd8112:data <=32'hFFBF00B6;14'd8113:data <=32'hFFE300BD;14'd8114:data <=32'h000400BB;
14'd8115:data <=32'h002300B2;14'd8116:data <=32'h003E00A4;14'd8117:data <=32'h00540091;
14'd8118:data <=32'h0065007B;14'd8119:data <=32'h006E0062;14'd8120:data <=32'h00710048;
14'd8121:data <=32'h006B0031;14'd8122:data <=32'h005E0020;14'd8123:data <=32'h004C0017;
14'd8124:data <=32'h003B0018;14'd8125:data <=32'h002E0023;14'd8126:data <=32'h002A0035;
14'd8127:data <=32'h00310049;14'd8128:data <=32'h0077005C;14'd8129:data <=32'h00960058;
14'd8130:data <=32'h00A1003E;14'd8131:data <=32'h00680024;14'd8132:data <=32'h009B0049;
14'd8133:data <=32'h00AD0032;14'd8134:data <=32'h00BB0017;14'd8135:data <=32'h00C0FFF9;
14'd8136:data <=32'h00C2FFD9;14'd8137:data <=32'h00BEFFBB;14'd8138:data <=32'h00B3FF9B;
14'd8139:data <=32'h00A2FF7D;14'd8140:data <=32'h0088FF63;14'd8141:data <=32'h0068FF4F;
14'd8142:data <=32'h0045FF46;14'd8143:data <=32'h0021FF46;14'd8144:data <=32'h0002FF50;
14'd8145:data <=32'hFFEAFF5F;14'd8146:data <=32'hFFDAFF6F;14'd8147:data <=32'hFFCFFF7F;
14'd8148:data <=32'hFFC8FF8C;14'd8149:data <=32'hFFC2FF95;14'd8150:data <=32'hFFBAFF9D;
14'd8151:data <=32'hFFB0FFA8;14'd8152:data <=32'hFFA7FFB4;14'd8153:data <=32'hFF9FFFC5;
14'd8154:data <=32'hFF9CFFD8;14'd8155:data <=32'hFF9FFFEB;14'd8156:data <=32'hFFA7FFFC;
14'd8157:data <=32'hFFB3000A;14'd8158:data <=32'hFFC10014;14'd8159:data <=32'hFFD00019;
14'd8160:data <=32'hFFE00019;14'd8161:data <=32'hFFEE0016;14'd8162:data <=32'hFFFD000F;
14'd8163:data <=32'h000A0004;14'd8164:data <=32'h0013FFF4;14'd8165:data <=32'h0017FFE0;
14'd8166:data <=32'h0014FFC8;14'd8167:data <=32'h0008FFAF;14'd8168:data <=32'hFFF1FF99;
14'd8169:data <=32'hFFD1FF8D;14'd8170:data <=32'hFFACFF8A;14'd8171:data <=32'hFF86FF95;
14'd8172:data <=32'hFF64FFAB;14'd8173:data <=32'hFF4AFFCD;14'd8174:data <=32'hFF3CFFF3;
14'd8175:data <=32'hFF39001C;14'd8176:data <=32'hFF3F0043;14'd8177:data <=32'hFF4E0065;
14'd8178:data <=32'hFF630081;14'd8179:data <=32'hFF7C0098;14'd8180:data <=32'hFF9900A9;
14'd8181:data <=32'hFFB600B3;14'd8182:data <=32'hFFD400B7;14'd8183:data <=32'hFFF100B5;
14'd8184:data <=32'h000C00AC;14'd8185:data <=32'h0020009E;14'd8186:data <=32'h002D008E;
14'd8187:data <=32'h0035007F;14'd8188:data <=32'h00360074;14'd8189:data <=32'h0036006F;
14'd8190:data <=32'h00370071;14'd8191:data <=32'h003F0076;14'd8192:data <=32'hFFF90039;
14'd8193:data <=32'hFFFD0059;14'd8194:data <=32'h0019006D;14'd8195:data <=32'h0084005D;
14'd8196:data <=32'h00B50075;14'd8197:data <=32'h00C20051;14'd8198:data <=32'h00C6002D;
14'd8199:data <=32'h00C0000A;14'd8200:data <=32'h00B4FFEE;14'd8201:data <=32'h00A4FFD7;
14'd8202:data <=32'h0093FFC5;14'd8203:data <=32'h0080FFB7;14'd8204:data <=32'h006CFFAD;
14'd8205:data <=32'h0057FFA8;14'd8206:data <=32'h0042FFAA;14'd8207:data <=32'h0032FFB1;
14'd8208:data <=32'h0027FFBD;14'd8209:data <=32'h0023FFCA;14'd8210:data <=32'h0028FFD5;
14'd8211:data <=32'h0032FFD9;14'd8212:data <=32'h003EFFD4;14'd8213:data <=32'h0046FFC8;
14'd8214:data <=32'h0048FFB5;14'd8215:data <=32'h0042FFA2;14'd8216:data <=32'h0033FF91;
14'd8217:data <=32'h001EFF87;14'd8218:data <=32'h0007FF83;14'd8219:data <=32'hFFEFFF87;
14'd8220:data <=32'hFFDCFF90;14'd8221:data <=32'hFFCDFF9E;14'd8222:data <=32'hFFC2FFAF;
14'd8223:data <=32'hFFBBFFC0;14'd8224:data <=32'hFFBAFFD3;14'd8225:data <=32'hFFBEFFE4;
14'd8226:data <=32'hFFC6FFF4;14'd8227:data <=32'hFFD30002;14'd8228:data <=32'hFFE50008;
14'd8229:data <=32'hFFF90007;14'd8230:data <=32'h000CFFFD;14'd8231:data <=32'h0019FFEC;
14'd8232:data <=32'h0020FFD6;14'd8233:data <=32'h001BFFBD;14'd8234:data <=32'h000EFFA8;
14'd8235:data <=32'hFFFAFF97;14'd8236:data <=32'hFFE2FF8F;14'd8237:data <=32'hFFC9FF8E;
14'd8238:data <=32'hFFB1FF94;14'd8239:data <=32'hFF9EFF9F;14'd8240:data <=32'hFF8EFFAB;
14'd8241:data <=32'hFF80FFB8;14'd8242:data <=32'hFF73FFC6;14'd8243:data <=32'hFF67FFD5;
14'd8244:data <=32'hFF5AFFE7;14'd8245:data <=32'hFF50FFFC;14'd8246:data <=32'hFF490015;
14'd8247:data <=32'hFF470030;14'd8248:data <=32'hFF4A004C;14'd8249:data <=32'hFF520067;
14'd8250:data <=32'hFF5D0080;14'd8251:data <=32'hFF6A0098;14'd8252:data <=32'hFF7A00B1;
14'd8253:data <=32'hFF8F00C9;14'd8254:data <=32'hFFAA00E2;14'd8255:data <=32'hFFCD00F7;
14'd8256:data <=32'hFFFD002C;14'd8257:data <=32'hFFEA0040;14'd8258:data <=32'hFFE40069;
14'd8259:data <=32'h002100FB;14'd8260:data <=32'h0076011A;14'd8261:data <=32'h00A700F3;
14'd8262:data <=32'h00C900C3;14'd8263:data <=32'h00DE008E;14'd8264:data <=32'h00E4005B;
14'd8265:data <=32'h00DE002C;14'd8266:data <=32'h00CF0004;14'd8267:data <=32'h00BAFFE2;
14'd8268:data <=32'h009FFFC7;14'd8269:data <=32'h007FFFB7;14'd8270:data <=32'h0060FFAE;
14'd8271:data <=32'h0040FFB1;14'd8272:data <=32'h0027FFBE;14'd8273:data <=32'h0016FFD1;
14'd8274:data <=32'h0010FFE7;14'd8275:data <=32'h0016FFFC;14'd8276:data <=32'h0023000A;
14'd8277:data <=32'h0035000D;14'd8278:data <=32'h00450008;14'd8279:data <=32'h0051FFFB;
14'd8280:data <=32'h0057FFEB;14'd8281:data <=32'h0056FFDB;14'd8282:data <=32'h0050FFCC;
14'd8283:data <=32'h0047FFC3;14'd8284:data <=32'h003EFFBA;14'd8285:data <=32'h0034FFB5;
14'd8286:data <=32'h002AFFB2;14'd8287:data <=32'h0021FFAF;14'd8288:data <=32'h0016FFAE;
14'd8289:data <=32'h000DFFB0;14'd8290:data <=32'h0002FFB3;14'd8291:data <=32'hFFFBFFBA;
14'd8292:data <=32'hFFF7FFC1;14'd8293:data <=32'hFFF7FFC8;14'd8294:data <=32'hFFF9FFCD;
14'd8295:data <=32'hFFFDFFCE;14'd8296:data <=32'h0000FFCC;14'd8297:data <=32'h0000FFC9;
14'd8298:data <=32'hFFFEFFC5;14'd8299:data <=32'hFFF9FFC1;14'd8300:data <=32'hFFF3FFC2;
14'd8301:data <=32'hFFF0FFC5;14'd8302:data <=32'hFFEFFFC8;14'd8303:data <=32'hFFF3FFC9;
14'd8304:data <=32'hFFF9FFC6;14'd8305:data <=32'hFFFDFFBC;14'd8306:data <=32'hFFFEFFAD;
14'd8307:data <=32'hFFF7FF9A;14'd8308:data <=32'hFFE8FF87;14'd8309:data <=32'hFFD1FF78;
14'd8310:data <=32'hFFB2FF6E;14'd8311:data <=32'hFF90FF6F;14'd8312:data <=32'hFF6BFF77;
14'd8313:data <=32'hFF48FF8A;14'd8314:data <=32'hFF27FFA3;14'd8315:data <=32'hFF0AFFC5;
14'd8316:data <=32'hFEF2FFF1;14'd8317:data <=32'hFEE40025;14'd8318:data <=32'hFEE1005E;
14'd8319:data <=32'hFEEE009C;14'd8320:data <=32'hFF93004E;14'd8321:data <=32'hFF860068;
14'd8322:data <=32'hFF72007E;14'd8323:data <=32'hFF3000C7;14'd8324:data <=32'hFF810118;
14'd8325:data <=32'hFFBC0120;14'd8326:data <=32'hFFF3011A;14'd8327:data <=32'h00250107;
14'd8328:data <=32'h004B00EE;14'd8329:data <=32'h006A00D1;14'd8330:data <=32'h008000B2;
14'd8331:data <=32'h00900092;14'd8332:data <=32'h009A0070;14'd8333:data <=32'h009B0050;
14'd8334:data <=32'h00960033;14'd8335:data <=32'h008A001A;14'd8336:data <=32'h007A0008;
14'd8337:data <=32'h0069FFFF;14'd8338:data <=32'h005CFFFB;14'd8339:data <=32'h0052FFFB;
14'd8340:data <=32'h004EFFFB;14'd8341:data <=32'h004DFFF9;14'd8342:data <=32'h004BFFF4;
14'd8343:data <=32'h0048FFEC;14'd8344:data <=32'h0041FFE4;14'd8345:data <=32'h0037FFE1;
14'd8346:data <=32'h002CFFE1;14'd8347:data <=32'h0022FFE7;14'd8348:data <=32'h001CFFEF;
14'd8349:data <=32'h001BFFFB;14'd8350:data <=32'h00210002;14'd8351:data <=32'h002A0007;
14'd8352:data <=32'h00340008;14'd8353:data <=32'h003E0004;14'd8354:data <=32'h0047FFFD;
14'd8355:data <=32'h004DFFF3;14'd8356:data <=32'h0051FFE8;14'd8357:data <=32'h0053FFDC;
14'd8358:data <=32'h0053FFCE;14'd8359:data <=32'h004FFFC0;14'd8360:data <=32'h0048FFB1;
14'd8361:data <=32'h003CFFA4;14'd8362:data <=32'h002BFF9B;14'd8363:data <=32'h0018FF97;
14'd8364:data <=32'h0004FF9A;14'd8365:data <=32'hFFF5FFA5;14'd8366:data <=32'hFFEBFFB4;
14'd8367:data <=32'hFFEBFFC5;14'd8368:data <=32'hFFF2FFD3;14'd8369:data <=32'h0000FFDB;
14'd8370:data <=32'h0011FFD7;14'd8371:data <=32'h001FFFCC;14'd8372:data <=32'h0028FFB8;
14'd8373:data <=32'h0028FFA0;14'd8374:data <=32'h001FFF88;14'd8375:data <=32'h000DFF71;
14'd8376:data <=32'hFFF4FF5D;14'd8377:data <=32'hFFD6FF51;14'd8378:data <=32'hFFB3FF4B;
14'd8379:data <=32'hFF8CFF4B;14'd8380:data <=32'hFF64FF57;14'd8381:data <=32'hFF3BFF6D;
14'd8382:data <=32'hFF17FF8E;14'd8383:data <=32'hFEFAFFBB;14'd8384:data <=32'hFF2CFFA4;
14'd8385:data <=32'hFEFEFFCA;14'd8386:data <=32'hFEECFFEB;14'd8387:data <=32'hFF16FFEC;
14'd8388:data <=32'hFF3A0044;14'd8389:data <=32'hFF4E005A;14'd8390:data <=32'hFF61006B;
14'd8391:data <=32'hFF740075;14'd8392:data <=32'hFF82007E;14'd8393:data <=32'hFF8F0089;
14'd8394:data <=32'hFF9D0096;14'd8395:data <=32'hFFAF00A3;14'd8396:data <=32'hFFC500AD;
14'd8397:data <=32'hFFDC00B4;14'd8398:data <=32'hFFF500B6;14'd8399:data <=32'h000E00B3;
14'd8400:data <=32'h002600AE;14'd8401:data <=32'h003B00A5;14'd8402:data <=32'h00510099;
14'd8403:data <=32'h0066008B;14'd8404:data <=32'h007A0077;14'd8405:data <=32'h008C005E;
14'd8406:data <=32'h0097003F;14'd8407:data <=32'h0099001C;14'd8408:data <=32'h008FFFF9;
14'd8409:data <=32'h007BFFDC;14'd8410:data <=32'h005FFFC9;14'd8411:data <=32'h003FFFC0;
14'd8412:data <=32'h0021FFC3;14'd8413:data <=32'h0008FFCF;14'd8414:data <=32'hFFF8FFE4;
14'd8415:data <=32'hFFF0FFF9;14'd8416:data <=32'hFFF1000F;14'd8417:data <=32'hFFF80022;
14'd8418:data <=32'h00040032;14'd8419:data <=32'h0014003C;14'd8420:data <=32'h00260042;
14'd8421:data <=32'h003A0043;14'd8422:data <=32'h004F003E;14'd8423:data <=32'h00630033;
14'd8424:data <=32'h00730021;14'd8425:data <=32'h007E000B;14'd8426:data <=32'h0081FFF3;
14'd8427:data <=32'h007DFFDC;14'd8428:data <=32'h0073FFC7;14'd8429:data <=32'h0065FFBA;
14'd8430:data <=32'h0056FFB3;14'd8431:data <=32'h004AFFB1;14'd8432:data <=32'h0044FFB1;
14'd8433:data <=32'h0041FFB1;14'd8434:data <=32'h0041FFAC;14'd8435:data <=32'h0043FFA4;
14'd8436:data <=32'h0041FF97;14'd8437:data <=32'h003BFF87;14'd8438:data <=32'h002EFF78;
14'd8439:data <=32'h001DFF6B;14'd8440:data <=32'h0009FF63;14'd8441:data <=32'hFFF3FF60;
14'd8442:data <=32'hFFDDFF5F;14'd8443:data <=32'hFFC8FF61;14'd8444:data <=32'hFFB2FF67;
14'd8445:data <=32'hFF9BFF6E;14'd8446:data <=32'hFF86FF7E;14'd8447:data <=32'hFF71FF90;
14'd8448:data <=32'hFFC1FF06;14'd8449:data <=32'hFF78FF01;14'd8450:data <=32'hFF41FF22;
14'd8451:data <=32'hFF79FFB4;14'd8452:data <=32'hFF99FFF6;14'd8453:data <=32'hFFA7FFF5;
14'd8454:data <=32'hFFAEFFED;14'd8455:data <=32'hFFAEFFE2;14'd8456:data <=32'hFFA4FFDA;
14'd8457:data <=32'hFF91FFD7;14'd8458:data <=32'hFF7CFFDE;14'd8459:data <=32'hFF68FFEF;
14'd8460:data <=32'hFF580008;14'd8461:data <=32'hFF510025;14'd8462:data <=32'hFF500045;
14'd8463:data <=32'hFF580065;14'd8464:data <=32'hFF670083;14'd8465:data <=32'hFF7D00A0;
14'd8466:data <=32'hFF9900B8;14'd8467:data <=32'hFFBD00CB;14'd8468:data <=32'hFFE600D5;
14'd8469:data <=32'h001300D4;14'd8470:data <=32'h003E00C5;14'd8471:data <=32'h006400AA;
14'd8472:data <=32'h007D0085;14'd8473:data <=32'h008B005C;14'd8474:data <=32'h008A0034;
14'd8475:data <=32'h007D0011;14'd8476:data <=32'h0069FFF7;14'd8477:data <=32'h0050FFE6;
14'd8478:data <=32'h0038FFE0;14'd8479:data <=32'h0022FFE0;14'd8480:data <=32'h000FFFE5;
14'd8481:data <=32'hFFFFFFEE;14'd8482:data <=32'hFFF3FFF9;14'd8483:data <=32'hFFEA0007;
14'd8484:data <=32'hFFE50017;14'd8485:data <=32'hFFE5002A;14'd8486:data <=32'hFFEB003C;
14'd8487:data <=32'hFFF6004D;14'd8488:data <=32'h0006005B;14'd8489:data <=32'h00190062;
14'd8490:data <=32'h002E0066;14'd8491:data <=32'h00430064;14'd8492:data <=32'h0056005E;
14'd8493:data <=32'h00670057;14'd8494:data <=32'h0079004D;14'd8495:data <=32'h008A0043;
14'd8496:data <=32'h009D0034;14'd8497:data <=32'h00B00021;14'd8498:data <=32'h00C20006;
14'd8499:data <=32'h00CFFFE3;14'd8500:data <=32'h00D3FFBB;14'd8501:data <=32'h00CBFF90;
14'd8502:data <=32'h00B7FF65;14'd8503:data <=32'h0099FF41;14'd8504:data <=32'h0071FF29;
14'd8505:data <=32'h0046FF19;14'd8506:data <=32'h001BFF15;14'd8507:data <=32'hFFF2FF1C;
14'd8508:data <=32'hFFCDFF29;14'd8509:data <=32'hFFADFF3D;14'd8510:data <=32'hFF92FF56;
14'd8511:data <=32'hFF7FFF75;14'd8512:data <=32'h004CFF4C;14'd8513:data <=32'h0025FF26;
14'd8514:data <=32'hFFE6FF18;14'd8515:data <=32'hFF77FF8B;14'd8516:data <=32'hFF98FFDD;
14'd8517:data <=32'hFFAEFFE7;14'd8518:data <=32'hFFC2FFE6;14'd8519:data <=32'hFFD1FFDD;
14'd8520:data <=32'hFFD6FFCD;14'd8521:data <=32'hFFCFFFBD;14'd8522:data <=32'hFFC1FFB3;
14'd8523:data <=32'hFFADFFAF;14'd8524:data <=32'hFF98FFB4;14'd8525:data <=32'hFF85FFBF;
14'd8526:data <=32'hFF74FFD0;14'd8527:data <=32'hFF68FFE4;14'd8528:data <=32'hFF60FFFB;
14'd8529:data <=32'hFF5C0015;14'd8530:data <=32'hFF5D0031;14'd8531:data <=32'hFF65004D;
14'd8532:data <=32'hFF740068;14'd8533:data <=32'hFF8C007F;14'd8534:data <=32'hFFAA008E;
14'd8535:data <=32'hFFCA0094;14'd8536:data <=32'hFFE80090;14'd8537:data <=32'h00020084;
14'd8538:data <=32'h00140075;14'd8539:data <=32'h001E0063;14'd8540:data <=32'h00230053;
14'd8541:data <=32'h00260047;14'd8542:data <=32'h0027003E;14'd8543:data <=32'h00280035;
14'd8544:data <=32'h002A002C;14'd8545:data <=32'h002A0021;14'd8546:data <=32'h00280016;
14'd8547:data <=32'h0020000A;14'd8548:data <=32'h00150001;14'd8549:data <=32'h0007FFFC;
14'd8550:data <=32'hFFF6FFFD;14'd8551:data <=32'hFFE70003;14'd8552:data <=32'hFFDA0010;
14'd8553:data <=32'hFFD00020;14'd8554:data <=32'hFFCB0033;14'd8555:data <=32'hFFCA0048;
14'd8556:data <=32'hFFCF005F;14'd8557:data <=32'hFFD90077;14'd8558:data <=32'hFFEB008F;
14'd8559:data <=32'h000400A6;14'd8560:data <=32'h002700B8;14'd8561:data <=32'h005200C1;
14'd8562:data <=32'h008300BD;14'd8563:data <=32'h00B400AB;14'd8564:data <=32'h00E20088;
14'd8565:data <=32'h0104005A;14'd8566:data <=32'h01190023;14'd8567:data <=32'h011EFFE6;
14'd8568:data <=32'h0113FFAD;14'd8569:data <=32'h00FAFF7A;14'd8570:data <=32'h00D8FF52;
14'd8571:data <=32'h00AFFF32;14'd8572:data <=32'h0083FF1D;14'd8573:data <=32'h0057FF13;
14'd8574:data <=32'h0029FF12;14'd8575:data <=32'hFFFFFF1A;14'd8576:data <=32'h0047FF71;
14'd8577:data <=32'h0036FF5B;14'd8578:data <=32'h001EFF3D;14'd8579:data <=32'hFFEDFF15;
14'd8580:data <=32'hFFEAFF5F;14'd8581:data <=32'hFFE1FF6B;14'd8582:data <=32'hFFDAFF72;
14'd8583:data <=32'hFFD4FF77;14'd8584:data <=32'hFFCBFF76;14'd8585:data <=32'hFFBCFF77;
14'd8586:data <=32'hFFA9FF7D;14'd8587:data <=32'hFF96FF89;14'd8588:data <=32'hFF85FF9B;
14'd8589:data <=32'hFF7AFFB0;14'd8590:data <=32'hFF75FFC9;14'd8591:data <=32'hFF76FFDE;
14'd8592:data <=32'hFF7BFFF1;14'd8593:data <=32'hFF830001;14'd8594:data <=32'hFF8B000F;
14'd8595:data <=32'hFF95001A;14'd8596:data <=32'hFF9F0024;14'd8597:data <=32'hFFAC002C;
14'd8598:data <=32'hFFB80030;14'd8599:data <=32'hFFC6002F;14'd8600:data <=32'hFFD0002A;
14'd8601:data <=32'hFFD70022;14'd8602:data <=32'hFFD6001A;14'd8603:data <=32'hFFD10014;
14'd8604:data <=32'hFFC80014;14'd8605:data <=32'hFFC2001B;14'd8606:data <=32'hFFBD0027;
14'd8607:data <=32'hFFBF0034;14'd8608:data <=32'hFFC80042;14'd8609:data <=32'hFFD50049;
14'd8610:data <=32'hFFE6004D;14'd8611:data <=32'hFFF50049;14'd8612:data <=32'h00020040;
14'd8613:data <=32'h00080033;14'd8614:data <=32'h00080026;14'd8615:data <=32'h0004001B;
14'd8616:data <=32'hFFFC0012;14'd8617:data <=32'hFFF0000D;14'd8618:data <=32'hFFE4000D;
14'd8619:data <=32'hFFD60011;14'd8620:data <=32'hFFC7001A;14'd8621:data <=32'hFFB90028;
14'd8622:data <=32'hFFB0003F;14'd8623:data <=32'hFFAC005A;14'd8624:data <=32'hFFB2007A;
14'd8625:data <=32'hFFC3009A;14'd8626:data <=32'hFFE100B6;14'd8627:data <=32'h000700C9;
14'd8628:data <=32'h003300D0;14'd8629:data <=32'h006000C9;14'd8630:data <=32'h008900B7;
14'd8631:data <=32'h00AA009C;14'd8632:data <=32'h00C2007B;14'd8633:data <=32'h00D10058;
14'd8634:data <=32'h00DA0037;14'd8635:data <=32'h00DE0016;14'd8636:data <=32'h00DDFFF7;
14'd8637:data <=32'h00D8FFDA;14'd8638:data <=32'h00CEFFBB;14'd8639:data <=32'h00C1FFA0;
14'd8640:data <=32'h00A6FF6D;14'd8641:data <=32'h0090FF51;14'd8642:data <=32'h0082FF48;
14'd8643:data <=32'h00C4FF7A;14'd8644:data <=32'h00C8FF99;14'd8645:data <=32'h00BFFF79;
14'd8646:data <=32'h00AFFF59;14'd8647:data <=32'h0099FF38;14'd8648:data <=32'h0078FF1A;
14'd8649:data <=32'h004DFF02;14'd8650:data <=32'h0019FEF5;14'd8651:data <=32'hFFE4FEF7;
14'd8652:data <=32'hFFB0FF09;14'd8653:data <=32'hFF84FF26;14'd8654:data <=32'hFF62FF4F;
14'd8655:data <=32'hFF50FF7C;14'd8656:data <=32'hFF4AFFA8;14'd8657:data <=32'hFF4EFFD0;
14'd8658:data <=32'hFF5BFFF3;14'd8659:data <=32'hFF6D000F;14'd8660:data <=32'hFF840026;
14'd8661:data <=32'hFF9F0035;14'd8662:data <=32'hFFBB003B;14'd8663:data <=32'hFFD70039;
14'd8664:data <=32'hFFF0002E;14'd8665:data <=32'h0001001B;14'd8666:data <=32'h00090004;
14'd8667:data <=32'h0007FFED;14'd8668:data <=32'hFFFAFFDA;14'd8669:data <=32'hFFE8FFD1;
14'd8670:data <=32'hFFD5FFCE;14'd8671:data <=32'hFFC2FFD5;14'd8672:data <=32'hFFB5FFE0;
14'd8673:data <=32'hFFAFFFEF;14'd8674:data <=32'hFFADFFFC;14'd8675:data <=32'hFFB00007;
14'd8676:data <=32'hFFB4000F;14'd8677:data <=32'hFFB70013;14'd8678:data <=32'hFFBA0017;
14'd8679:data <=32'hFFBA001B;14'd8680:data <=32'hFFBA0020;14'd8681:data <=32'hFFBB0025;
14'd8682:data <=32'hFFBC0029;14'd8683:data <=32'hFFBD002E;14'd8684:data <=32'hFFBF0033;
14'd8685:data <=32'hFFBE0038;14'd8686:data <=32'hFFBE003E;14'd8687:data <=32'hFFBD0048;
14'd8688:data <=32'hFFBE0054;14'd8689:data <=32'hFFC30063;14'd8690:data <=32'hFFCC0072;
14'd8691:data <=32'hFFDC007E;14'd8692:data <=32'hFFEE0084;14'd8693:data <=32'h00020086;
14'd8694:data <=32'h00140082;14'd8695:data <=32'h0020007A;14'd8696:data <=32'h00280073;
14'd8697:data <=32'h002C006F;14'd8698:data <=32'h002E006F;14'd8699:data <=32'h00340074;
14'd8700:data <=32'h003F007B;14'd8701:data <=32'h00500082;14'd8702:data <=32'h00660084;
14'd8703:data <=32'h0080007F;14'd8704:data <=32'h00E80021;14'd8705:data <=32'h00F0FFFC;
14'd8706:data <=32'h00DEFFEA;14'd8707:data <=32'h00A8005B;14'd8708:data <=32'h00D4007F;
14'd8709:data <=32'h00F6005D;14'd8710:data <=32'h01120030;14'd8711:data <=32'h0123FFFB;
14'd8712:data <=32'h0125FFBF;14'd8713:data <=32'h0116FF81;14'd8714:data <=32'h00F6FF47;
14'd8715:data <=32'h00C7FF1A;14'd8716:data <=32'h008DFEFC;14'd8717:data <=32'h0051FEF0;
14'd8718:data <=32'h0017FEF5;14'd8719:data <=32'hFFE4FF07;14'd8720:data <=32'hFFBBFF21;
14'd8721:data <=32'hFF9BFF42;14'd8722:data <=32'hFF86FF65;14'd8723:data <=32'hFF79FF88;
14'd8724:data <=32'hFF74FFAD;14'd8725:data <=32'hFF78FFCF;14'd8726:data <=32'hFF84FFEF;
14'd8727:data <=32'hFF970007;14'd8728:data <=32'hFFAF0018;14'd8729:data <=32'hFFC9001E;
14'd8730:data <=32'hFFE0001C;14'd8731:data <=32'hFFF20013;14'd8732:data <=32'hFFFE0006;
14'd8733:data <=32'h0002FFF8;14'd8734:data <=32'h0003FFED;14'd8735:data <=32'h0000FFE5;
14'd8736:data <=32'hFFFEFFDE;14'd8737:data <=32'hFFFCFFD8;14'd8738:data <=32'hFFFAFFD1;
14'd8739:data <=32'hFFF6FFC9;14'd8740:data <=32'hFFEFFFBD;14'd8741:data <=32'hFFE3FFB3;
14'd8742:data <=32'hFFD2FFAC;14'd8743:data <=32'hFFBDFFAA;14'd8744:data <=32'hFFA6FFAD;
14'd8745:data <=32'hFF91FFB9;14'd8746:data <=32'hFF7EFFCA;14'd8747:data <=32'hFF6FFFE0;
14'd8748:data <=32'hFF67FFF9;14'd8749:data <=32'hFF640013;14'd8750:data <=32'hFF66002C;
14'd8751:data <=32'hFF6E0045;14'd8752:data <=32'hFF7A005C;14'd8753:data <=32'hFF8B0071;
14'd8754:data <=32'hFFA10083;14'd8755:data <=32'hFFBB008E;14'd8756:data <=32'hFFD90090;
14'd8757:data <=32'hFFF30089;14'd8758:data <=32'h0009007A;14'd8759:data <=32'h00150066;
14'd8760:data <=32'h00180051;14'd8761:data <=32'h000F0040;14'd8762:data <=32'h00010039;
14'd8763:data <=32'hFFF1003A;14'd8764:data <=32'hFFE20047;14'd8765:data <=32'hFFDC005B;
14'd8766:data <=32'hFFDF0073;14'd8767:data <=32'hFFEB008B;14'd8768:data <=32'h0039009F;
14'd8769:data <=32'h005200A6;14'd8770:data <=32'h005E0095;14'd8771:data <=32'h00230078;
14'd8772:data <=32'h004800B9;14'd8773:data <=32'h006C00B7;14'd8774:data <=32'h009200AA;
14'd8775:data <=32'h00B50094;14'd8776:data <=32'h00D30070;14'd8777:data <=32'h00E90045;
14'd8778:data <=32'h00F10017;14'd8779:data <=32'h00EAFFE9;14'd8780:data <=32'h00D9FFC0;
14'd8781:data <=32'h00C0FF9F;14'd8782:data <=32'h00A4FF8A;14'd8783:data <=32'h0087FF7D;
14'd8784:data <=32'h006FFF75;14'd8785:data <=32'h0058FF71;14'd8786:data <=32'h0041FF6E;
14'd8787:data <=32'h002DFF6D;14'd8788:data <=32'h0016FF6F;14'd8789:data <=32'h0001FF75;
14'd8790:data <=32'hFFEFFF80;14'd8791:data <=32'hFFDFFF8D;14'd8792:data <=32'hFFD4FF9C;
14'd8793:data <=32'hFFCEFFAC;14'd8794:data <=32'hFFCBFFBA;14'd8795:data <=32'hFFC9FFC6;
14'd8796:data <=32'hFFC9FFD2;14'd8797:data <=32'hFFC9FFDE;14'd8798:data <=32'hFFCCFFEC;
14'd8799:data <=32'hFFD3FFF9;14'd8800:data <=32'hFFDF0006;14'd8801:data <=32'hFFF0000E;
14'd8802:data <=32'h0006000F;14'd8803:data <=32'h001B0007;14'd8804:data <=32'h002FFFF7;
14'd8805:data <=32'h003BFFDD;14'd8806:data <=32'h003CFFC0;14'd8807:data <=32'h0034FFA1;
14'd8808:data <=32'h0021FF87;14'd8809:data <=32'h0005FF73;14'd8810:data <=32'hFFE4FF69;
14'd8811:data <=32'hFFC3FF67;14'd8812:data <=32'hFFA2FF6F;14'd8813:data <=32'hFF84FF7E;
14'd8814:data <=32'hFF69FF93;14'd8815:data <=32'hFF53FFAF;14'd8816:data <=32'hFF43FFCE;
14'd8817:data <=32'hFF3CFFF2;14'd8818:data <=32'hFF3E0017;14'd8819:data <=32'hFF490039;
14'd8820:data <=32'hFF5D0055;14'd8821:data <=32'hFF76006A;14'd8822:data <=32'hFF930074;
14'd8823:data <=32'hFFAC0075;14'd8824:data <=32'hFFBE006E;14'd8825:data <=32'hFFC90064;
14'd8826:data <=32'hFFCD005D;14'd8827:data <=32'hFFCA005A;14'd8828:data <=32'hFFC7005E;
14'd8829:data <=32'hFFC60068;14'd8830:data <=32'hFFC90076;14'd8831:data <=32'hFFD10084;
14'd8832:data <=32'hFFB70035;14'd8833:data <=32'hFFAB0055;14'd8834:data <=32'hFFB6006F;
14'd8835:data <=32'h0013007F;14'd8836:data <=32'h002E00B5;14'd8837:data <=32'h004600AB;
14'd8838:data <=32'h005E009D;14'd8839:data <=32'h0072008B;14'd8840:data <=32'h00820074;
14'd8841:data <=32'h008E0058;14'd8842:data <=32'h008F003C;14'd8843:data <=32'h00890023;
14'd8844:data <=32'h007C000E;14'd8845:data <=32'h006C0004;14'd8846:data <=32'h005E0001;
14'd8847:data <=32'h00550005;14'd8848:data <=32'h0054000B;14'd8849:data <=32'h0058000E;
14'd8850:data <=32'h0062000D;14'd8851:data <=32'h006C0005;14'd8852:data <=32'h0074FFF7;
14'd8853:data <=32'h0077FFE6;14'd8854:data <=32'h0076FFD3;14'd8855:data <=32'h0070FFC1;
14'd8856:data <=32'h0066FFB1;14'd8857:data <=32'h0058FFA3;14'd8858:data <=32'h0048FF97;
14'd8859:data <=32'h0035FF8E;14'd8860:data <=32'h001DFF8A;14'd8861:data <=32'h0006FF8C;
14'd8862:data <=32'hFFEEFF96;14'd8863:data <=32'hFFDAFFA7;14'd8864:data <=32'hFFCDFFBF;
14'd8865:data <=32'hFFCBFFD9;14'd8866:data <=32'hFFD3FFF2;14'd8867:data <=32'hFFE30007;
14'd8868:data <=32'hFFFB0010;14'd8869:data <=32'h00140011;14'd8870:data <=32'h002B0007;
14'd8871:data <=32'h003CFFF7;14'd8872:data <=32'h0047FFE0;14'd8873:data <=32'h0048FFC9;
14'd8874:data <=32'h0044FFB2;14'd8875:data <=32'h003AFF9E;14'd8876:data <=32'h002DFF8C;
14'd8877:data <=32'h001BFF7D;14'd8878:data <=32'h0007FF71;14'd8879:data <=32'hFFF0FF69;
14'd8880:data <=32'hFFD6FF65;14'd8881:data <=32'hFFBCFF67;14'd8882:data <=32'hFFA2FF70;
14'd8883:data <=32'hFF8AFF7E;14'd8884:data <=32'hFF76FF90;14'd8885:data <=32'hFF69FFA3;
14'd8886:data <=32'hFF5FFFB5;14'd8887:data <=32'hFF55FFC7;14'd8888:data <=32'hFF4EFFD7;
14'd8889:data <=32'hFF44FFEA;14'd8890:data <=32'hFF370000;14'd8891:data <=32'hFF2E001B;
14'd8892:data <=32'hFF29003D;14'd8893:data <=32'hFF2C0063;14'd8894:data <=32'hFF3B008B;
14'd8895:data <=32'hFF5400AF;14'd8896:data <=32'hFFD30000;14'd8897:data <=32'hFFB10006;
14'd8898:data <=32'hFF930025;14'd8899:data <=32'hFF9B00C6;14'd8900:data <=32'hFFCD0108;
14'd8901:data <=32'hFFFF0102;14'd8902:data <=32'h002E00F1;14'd8903:data <=32'h005300D7;
14'd8904:data <=32'h007300B6;14'd8905:data <=32'h0088008F;14'd8906:data <=32'h00910066;
14'd8907:data <=32'h008C003D;14'd8908:data <=32'h007C001C;14'd8909:data <=32'h00630005;
14'd8910:data <=32'h0047FFFC;14'd8911:data <=32'h002E0000;14'd8912:data <=32'h001D000C;
14'd8913:data <=32'h0016001C;14'd8914:data <=32'h0018002D;14'd8915:data <=32'h00220038;
14'd8916:data <=32'h0031003E;14'd8917:data <=32'h0040003F;14'd8918:data <=32'h004E0039;
14'd8919:data <=32'h005B0031;14'd8920:data <=32'h00650026;14'd8921:data <=32'h006D0017;
14'd8922:data <=32'h00730006;14'd8923:data <=32'h0075FFF3;14'd8924:data <=32'h0070FFDF;
14'd8925:data <=32'h0066FFCC;14'd8926:data <=32'h0056FFBE;14'd8927:data <=32'h0043FFB6;
14'd8928:data <=32'h0030FFB5;14'd8929:data <=32'h001FFFBA;14'd8930:data <=32'h0014FFC5;
14'd8931:data <=32'h000EFFD1;14'd8932:data <=32'h000EFFDC;14'd8933:data <=32'h0013FFE3;
14'd8934:data <=32'h0019FFE5;14'd8935:data <=32'h001EFFE4;14'd8936:data <=32'h0020FFE2;
14'd8937:data <=32'h0020FFE0;14'd8938:data <=32'h0020FFE0;14'd8939:data <=32'h0022FFE0;
14'd8940:data <=32'h0026FFE0;14'd8941:data <=32'h002DFFE0;14'd8942:data <=32'h0036FFDB;
14'd8943:data <=32'h003FFFD2;14'd8944:data <=32'h0046FFC3;14'd8945:data <=32'h0049FFB1;
14'd8946:data <=32'h0048FF9C;14'd8947:data <=32'h0041FF87;14'd8948:data <=32'h0035FF70;
14'd8949:data <=32'h0025FF5C;14'd8950:data <=32'h000FFF47;14'd8951:data <=32'hFFF3FF35;
14'd8952:data <=32'hFFCFFF27;14'd8953:data <=32'hFFA4FF1F;14'd8954:data <=32'hFF73FF22;
14'd8955:data <=32'hFF3EFF33;14'd8956:data <=32'hFF0CFF54;14'd8957:data <=32'hFEE2FF84;
14'd8958:data <=32'hFEC5FFC1;14'd8959:data <=32'hFEBC0004;14'd8960:data <=32'hFF8FFFF9;
14'd8961:data <=32'hFF79FFFE;14'd8962:data <=32'hFF540001;14'd8963:data <=32'hFEEB0035;
14'd8964:data <=32'hFF0A009E;14'd8965:data <=32'hFF3300C1;14'd8966:data <=32'hFF6100D9;
14'd8967:data <=32'hFF8F00E6;14'd8968:data <=32'hFFC000E8;14'd8969:data <=32'hFFED00DF;
14'd8970:data <=32'h001400CA;14'd8971:data <=32'h003000AF;14'd8972:data <=32'h00410090;
14'd8973:data <=32'h00470073;14'd8974:data <=32'h0043005C;14'd8975:data <=32'h003C004D;
14'd8976:data <=32'h00350045;14'd8977:data <=32'h00310041;14'd8978:data <=32'h00300041;
14'd8979:data <=32'h0034003E;14'd8980:data <=32'h0037003A;14'd8981:data <=32'h003A0033;
14'd8982:data <=32'h003A002B;14'd8983:data <=32'h00380025;14'd8984:data <=32'h00350020;
14'd8985:data <=32'h0032001E;14'd8986:data <=32'h0030001E;14'd8987:data <=32'h0030001D;
14'd8988:data <=32'h0032001D;14'd8989:data <=32'h0034001B;14'd8990:data <=32'h00350019;
14'd8991:data <=32'h00350017;14'd8992:data <=32'h00350018;14'd8993:data <=32'h00370018;
14'd8994:data <=32'h003C001A;14'd8995:data <=32'h0043001A;14'd8996:data <=32'h004D0016;
14'd8997:data <=32'h0057000D;14'd8998:data <=32'h005DFFFF;14'd8999:data <=32'h005FFFEE;
14'd9000:data <=32'h005AFFDD;14'd9001:data <=32'h004FFFCF;14'd9002:data <=32'h0040FFC7;
14'd9003:data <=32'h002FFFC6;14'd9004:data <=32'h0021FFCD;14'd9005:data <=32'h0019FFD9;
14'd9006:data <=32'h0018FFE6;14'd9007:data <=32'h001FFFF1;14'd9008:data <=32'h002BFFF9;
14'd9009:data <=32'h003AFFFB;14'd9010:data <=32'h004BFFF7;14'd9011:data <=32'h005CFFED;
14'd9012:data <=32'h006BFFDD;14'd9013:data <=32'h0077FFC5;14'd9014:data <=32'h007FFFA9;
14'd9015:data <=32'h0080FF87;14'd9016:data <=32'h0076FF60;14'd9017:data <=32'h0060FF39;
14'd9018:data <=32'h003DFF15;14'd9019:data <=32'h000EFEFC;14'd9020:data <=32'hFFD5FEF0;
14'd9021:data <=32'hFF9AFEF5;14'd9022:data <=32'hFF62FF0B;14'd9023:data <=32'hFF32FF2E;
14'd9024:data <=32'hFF7AFF4D;14'd9025:data <=32'hFF4AFF56;14'd9026:data <=32'hFF30FF5D;
14'd9027:data <=32'hFF41FF58;14'd9028:data <=32'hFF33FFB3;14'd9029:data <=32'hFF2FFFD0;
14'd9030:data <=32'hFF2EFFEE;14'd9031:data <=32'hFF310008;14'd9032:data <=32'hFF390024;
14'd9033:data <=32'hFF45003D;14'd9034:data <=32'hFF550052;14'd9035:data <=32'hFF660062;
14'd9036:data <=32'hFF76006E;14'd9037:data <=32'hFF84007A;14'd9038:data <=32'hFF920085;
14'd9039:data <=32'hFFA00093;14'd9040:data <=32'hFFB4009F;14'd9041:data <=32'hFFCD00AB;
14'd9042:data <=32'hFFEB00B2;14'd9043:data <=32'h000C00B0;14'd9044:data <=32'h002C00A4;
14'd9045:data <=32'h0048008E;14'd9046:data <=32'h005C0072;14'd9047:data <=32'h00650053;
14'd9048:data <=32'h00630036;14'd9049:data <=32'h005A001B;14'd9050:data <=32'h004C0008;
14'd9051:data <=32'h003AFFFC;14'd9052:data <=32'h0028FFF4;14'd9053:data <=32'h0016FFF3;
14'd9054:data <=32'h0005FFF7;14'd9055:data <=32'hFFF70000;14'd9056:data <=32'hFFEA000F;
14'd9057:data <=32'hFFE40022;14'd9058:data <=32'hFFE60037;14'd9059:data <=32'hFFF0004C;
14'd9060:data <=32'h0001005B;14'd9061:data <=32'h00180065;14'd9062:data <=32'h00330065;
14'd9063:data <=32'h004A005B;14'd9064:data <=32'h005C004C;14'd9065:data <=32'h00670038;
14'd9066:data <=32'h006A0024;14'd9067:data <=32'h00680014;14'd9068:data <=32'h00620009;
14'd9069:data <=32'h005C0004;14'd9070:data <=32'h00570000;14'd9071:data <=32'h0057FFFF;
14'd9072:data <=32'h0059FFFE;14'd9073:data <=32'h005DFFFA;14'd9074:data <=32'h0063FFF5;
14'd9075:data <=32'h0068FFED;14'd9076:data <=32'h006DFFE5;14'd9077:data <=32'h0072FFD9;
14'd9078:data <=32'h0076FFCD;14'd9079:data <=32'h007AFFBB;14'd9080:data <=32'h007BFFA6;
14'd9081:data <=32'h0078FF8E;14'd9082:data <=32'h006CFF73;14'd9083:data <=32'h0056FF5A;
14'd9084:data <=32'h003BFF49;14'd9085:data <=32'h0019FF3E;14'd9086:data <=32'hFFF9FF3F;
14'd9087:data <=32'hFFDAFF47;14'd9088:data <=32'h0044FEFC;14'd9089:data <=32'h000DFED9;
14'd9090:data <=32'hFFDBFEDA;14'd9091:data <=32'hFFE5FF5E;14'd9092:data <=32'hFFDDFF9A;
14'd9093:data <=32'hFFDDFF93;14'd9094:data <=32'hFFD5FF8C;14'd9095:data <=32'hFFC9FF84;
14'd9096:data <=32'hFFB6FF81;14'd9097:data <=32'hFFA2FF80;14'd9098:data <=32'hFF8DFF85;
14'd9099:data <=32'hFF75FF8E;14'd9100:data <=32'hFF5DFF9D;14'd9101:data <=32'hFF45FFB1;
14'd9102:data <=32'hFF30FFCE;14'd9103:data <=32'hFF20FFF3;14'd9104:data <=32'hFF1A001F;
14'd9105:data <=32'hFF20004E;14'd9106:data <=32'hFF35007C;14'd9107:data <=32'hFF5700A2;
14'd9108:data <=32'hFF8300BC;14'd9109:data <=32'hFFB300C7;14'd9110:data <=32'hFFE200C4;
14'd9111:data <=32'h000B00B5;14'd9112:data <=32'h002B009D;14'd9113:data <=32'h00400080;
14'd9114:data <=32'h004E0062;14'd9115:data <=32'h00530044;14'd9116:data <=32'h004F0029;
14'd9117:data <=32'h00470010;14'd9118:data <=32'h0039FFFC;14'd9119:data <=32'h0025FFEE;
14'd9120:data <=32'h000DFFE6;14'd9121:data <=32'hFFF5FFE7;14'd9122:data <=32'hFFDFFFF0;
14'd9123:data <=32'hFFCE0000;14'd9124:data <=32'hFFC40015;14'd9125:data <=32'hFFC2002C;
14'd9126:data <=32'hFFC70041;14'd9127:data <=32'hFFD20051;14'd9128:data <=32'hFFDE005D;
14'd9129:data <=32'hFFEB0065;14'd9130:data <=32'hFFF7006D;14'd9131:data <=32'h00020074;
14'd9132:data <=32'h000F007B;14'd9133:data <=32'h00210082;14'd9134:data <=32'h00340089;
14'd9135:data <=32'h004E008C;14'd9136:data <=32'h006A0087;14'd9137:data <=32'h0087007A;
14'd9138:data <=32'h00A10067;14'd9139:data <=32'h00B7004C;14'd9140:data <=32'h00C6002C;
14'd9141:data <=32'h00CD000B;14'd9142:data <=32'h00CEFFE9;14'd9143:data <=32'h00C9FFC9;
14'd9144:data <=32'h00BDFFA9;14'd9145:data <=32'h00ACFF8A;14'd9146:data <=32'h0095FF70;
14'd9147:data <=32'h0077FF5C;14'd9148:data <=32'h0054FF4F;14'd9149:data <=32'h002FFF4E;
14'd9150:data <=32'h000CFF57;14'd9151:data <=32'hFFF1FF6A;14'd9152:data <=32'h00B4FF8E;
14'd9153:data <=32'h00ACFF5B;14'd9154:data <=32'h0082FF33;14'd9155:data <=32'hFFFAFF7A;
14'd9156:data <=32'hFFFCFFC0;14'd9157:data <=32'h000BFFC2;14'd9158:data <=32'h0016FFBB;
14'd9159:data <=32'h001CFFAC;14'd9160:data <=32'h001BFF9D;14'd9161:data <=32'h0016FF8C;
14'd9162:data <=32'h0009FF7D;14'd9163:data <=32'hFFF8FF70;14'd9164:data <=32'hFFE1FF64;
14'd9165:data <=32'hFFC5FF5D;14'd9166:data <=32'hFFA4FF5E;14'd9167:data <=32'hFF82FF69;
14'd9168:data <=32'hFF60FF80;14'd9169:data <=32'hFF46FFA1;14'd9170:data <=32'hFF37FFC9;
14'd9171:data <=32'hFF34FFF4;14'd9172:data <=32'hFF3E001C;14'd9173:data <=32'hFF53003D;
14'd9174:data <=32'hFF6C0055;14'd9175:data <=32'hFF870063;14'd9176:data <=32'hFFA2006B;
14'd9177:data <=32'hFFB9006C;14'd9178:data <=32'hFFCD006B;14'd9179:data <=32'hFFE00067;
14'd9180:data <=32'hFFF10060;14'd9181:data <=32'h00020057;14'd9182:data <=32'h000E004A;
14'd9183:data <=32'h0017003A;14'd9184:data <=32'h001A0029;14'd9185:data <=32'h00190019;
14'd9186:data <=32'h0012000A;14'd9187:data <=32'h00080000;14'd9188:data <=32'hFFFCFFF9;
14'd9189:data <=32'hFFEFFFF6;14'd9190:data <=32'hFFE3FFF5;14'd9191:data <=32'hFFD6FFF6;
14'd9192:data <=32'hFFC8FFFA;14'd9193:data <=32'hFFB80000;14'd9194:data <=32'hFFA7000C;
14'd9195:data <=32'hFF980020;14'd9196:data <=32'hFF8C003B;14'd9197:data <=32'hFF86005D;
14'd9198:data <=32'hFF8D0085;14'd9199:data <=32'hFFA100AB;14'd9200:data <=32'hFFC200CC;
14'd9201:data <=32'hFFEB00E5;14'd9202:data <=32'h001D00F1;14'd9203:data <=32'h005000EF;
14'd9204:data <=32'h008100E0;14'd9205:data <=32'h00AD00C7;14'd9206:data <=32'h00D200A3;
14'd9207:data <=32'h00EE007A;14'd9208:data <=32'h0100004B;14'd9209:data <=32'h0108001A;
14'd9210:data <=32'h0105FFE8;14'd9211:data <=32'h00F4FFB8;14'd9212:data <=32'h00D8FF8E;
14'd9213:data <=32'h00B3FF6F;14'd9214:data <=32'h0089FF5D;14'd9215:data <=32'h005EFF5B;
14'd9216:data <=32'h0081FFD1;14'd9217:data <=32'h0089FFBE;14'd9218:data <=32'h008BFF9A;
14'd9219:data <=32'h0068FF5B;14'd9220:data <=32'h0053FF97;14'd9221:data <=32'h004FFF94;
14'd9222:data <=32'h0048FF8E;14'd9223:data <=32'h0040FF84;14'd9224:data <=32'h0033FF7C;
14'd9225:data <=32'h0025FF76;14'd9226:data <=32'h0015FF74;14'd9227:data <=32'h0006FF73;
14'd9228:data <=32'hFFF7FF73;14'd9229:data <=32'hFFE7FF74;14'd9230:data <=32'hFFD7FF77;
14'd9231:data <=32'hFFC5FF7D;14'd9232:data <=32'hFFB2FF89;14'd9233:data <=32'hFFA2FF99;
14'd9234:data <=32'hFF97FFAE;14'd9235:data <=32'hFF95FFC4;14'd9236:data <=32'hFF98FFD8;
14'd9237:data <=32'hFFA2FFE6;14'd9238:data <=32'hFFACFFEF;14'd9239:data <=32'hFFB6FFF2;
14'd9240:data <=32'hFFBBFFF0;14'd9241:data <=32'hFFBCFFEF;14'd9242:data <=32'hFFB7FFEF;
14'd9243:data <=32'hFFB1FFF3;14'd9244:data <=32'hFFADFFFC;14'd9245:data <=32'hFFAC0007;
14'd9246:data <=32'hFFAF0014;14'd9247:data <=32'hFFB5001D;14'd9248:data <=32'hFFBE0025;
14'd9249:data <=32'hFFC9002A;14'd9250:data <=32'hFFD3002C;14'd9251:data <=32'hFFDD002A;
14'd9252:data <=32'hFFE80027;14'd9253:data <=32'hFFF10022;14'd9254:data <=32'hFFF70017;
14'd9255:data <=32'hFFFB000A;14'd9256:data <=32'hFFF9FFFA;14'd9257:data <=32'hFFF0FFEA;
14'd9258:data <=32'hFFE0FFDD;14'd9259:data <=32'hFFC6FFD5;14'd9260:data <=32'hFFA9FFD8;
14'd9261:data <=32'hFF8BFFE6;14'd9262:data <=32'hFF710000;14'd9263:data <=32'hFF610025;
14'd9264:data <=32'hFF5D004E;14'd9265:data <=32'hFF650077;14'd9266:data <=32'hFF79009C;
14'd9267:data <=32'hFF9700BC;14'd9268:data <=32'hFFB900D4;14'd9269:data <=32'hFFE000E1;
14'd9270:data <=32'h000800E7;14'd9271:data <=32'h002F00E6;14'd9272:data <=32'h005600DD;
14'd9273:data <=32'h007B00CC;14'd9274:data <=32'h009B00B4;14'd9275:data <=32'h00B50095;
14'd9276:data <=32'h00C60072;14'd9277:data <=32'h00CE004F;14'd9278:data <=32'h00CD002D;
14'd9279:data <=32'h00C60012;14'd9280:data <=32'h00ADFFDF;14'd9281:data <=32'h00A5FFCF;
14'd9282:data <=32'h00AAFFCD;14'd9283:data <=32'h00E70007;14'd9284:data <=32'h00E80023;
14'd9285:data <=32'h00F5FFFD;14'd9286:data <=32'h00F7FFD2;14'd9287:data <=32'h00EFFFA4;
14'd9288:data <=32'h00D9FF79;14'd9289:data <=32'h00B9FF55;14'd9290:data <=32'h0092FF3B;
14'd9291:data <=32'h0069FF2C;14'd9292:data <=32'h003EFF27;14'd9293:data <=32'h0016FF2A;
14'd9294:data <=32'hFFF0FF35;14'd9295:data <=32'hFFCEFF47;14'd9296:data <=32'hFFB2FF5F;
14'd9297:data <=32'hFF9CFF7E;14'd9298:data <=32'hFF92FFA1;14'd9299:data <=32'hFF92FFC5;
14'd9300:data <=32'hFF9DFFE5;14'd9301:data <=32'hFFB1FFFC;14'd9302:data <=32'hFFCC0009;
14'd9303:data <=32'hFFE60009;14'd9304:data <=32'hFFF9FFFF;14'd9305:data <=32'h0006FFEF;
14'd9306:data <=32'h0009FFDE;14'd9307:data <=32'h0004FFCE;14'd9308:data <=32'hFFFAFFC2;
14'd9309:data <=32'hFFEDFFBD;14'd9310:data <=32'hFFE0FFBC;14'd9311:data <=32'hFFD4FFBF;
14'd9312:data <=32'hFFCBFFC5;14'd9313:data <=32'hFFC2FFCA;14'd9314:data <=32'hFFBCFFD3;
14'd9315:data <=32'hFFB8FFDC;14'd9316:data <=32'hFFB5FFE7;14'd9317:data <=32'hFFB7FFF1;
14'd9318:data <=32'hFFBBFFF9;14'd9319:data <=32'hFFC1FFFE;14'd9320:data <=32'hFFCAFFFE;
14'd9321:data <=32'hFFCEFFFB;14'd9322:data <=32'hFFD0FFF4;14'd9323:data <=32'hFFCBFFEB;
14'd9324:data <=32'hFFC0FFE7;14'd9325:data <=32'hFFB2FFE6;14'd9326:data <=32'hFFA2FFED;
14'd9327:data <=32'hFF95FFFA;14'd9328:data <=32'hFF8B000C;14'd9329:data <=32'hFF88001F;
14'd9330:data <=32'hFF8C0032;14'd9331:data <=32'hFF920042;14'd9332:data <=32'hFF9A004F;
14'd9333:data <=32'hFFA10058;14'd9334:data <=32'hFFA70062;14'd9335:data <=32'hFFAD006C;
14'd9336:data <=32'hFFB30078;14'd9337:data <=32'hFFBB0085;14'd9338:data <=32'hFFC70093;
14'd9339:data <=32'hFFD600A0;14'd9340:data <=32'hFFE700AB;14'd9341:data <=32'hFFFA00B3;
14'd9342:data <=32'h000D00BB;14'd9343:data <=32'h002400C2;14'd9344:data <=32'h00A0007A;
14'd9345:data <=32'h00AC0069;14'd9346:data <=32'h00A40063;14'd9347:data <=32'h005B00CD;
14'd9348:data <=32'h00810102;14'd9349:data <=32'h00BA00EC;14'd9350:data <=32'h00ED00C6;
14'd9351:data <=32'h01160092;14'd9352:data <=32'h012D0056;14'd9353:data <=32'h01340016;
14'd9354:data <=32'h0129FFD9;14'd9355:data <=32'h0113FFA3;14'd9356:data <=32'h00F3FF76;
14'd9357:data <=32'h00CAFF53;14'd9358:data <=32'h009EFF39;14'd9359:data <=32'h006DFF2B;
14'd9360:data <=32'h003CFF29;14'd9361:data <=32'h000DFF33;14'd9362:data <=32'hFFE4FF48;
14'd9363:data <=32'hFFC6FF67;14'd9364:data <=32'hFFB3FF8B;14'd9365:data <=32'hFFAFFFB0;
14'd9366:data <=32'hFFB6FFCF;14'd9367:data <=32'hFFC5FFE7;14'd9368:data <=32'hFFD7FFF4;
14'd9369:data <=32'hFFE8FFF9;14'd9370:data <=32'hFFF7FFF9;14'd9371:data <=32'h0001FFF5;
14'd9372:data <=32'h0008FFF0;14'd9373:data <=32'h000CFFEB;14'd9374:data <=32'h0011FFE6;
14'd9375:data <=32'h0016FFE0;14'd9376:data <=32'h0019FFD9;14'd9377:data <=32'h001BFFCF;
14'd9378:data <=32'h0019FFC3;14'd9379:data <=32'h0014FFB7;14'd9380:data <=32'h000CFFAC;
14'd9381:data <=32'h0000FFA5;14'd9382:data <=32'hFFF3FF9F;14'd9383:data <=32'hFFE5FF9D;
14'd9384:data <=32'hFFD8FF9C;14'd9385:data <=32'hFFCAFF9D;14'd9386:data <=32'hFFBAFF9F;
14'd9387:data <=32'hFFAAFFA4;14'd9388:data <=32'hFF99FFAD;14'd9389:data <=32'hFF89FFBA;
14'd9390:data <=32'hFF7AFFCD;14'd9391:data <=32'hFF70FFE6;14'd9392:data <=32'hFF700000;
14'd9393:data <=32'hFF78001A;14'd9394:data <=32'hFF87002E;14'd9395:data <=32'hFF9A003B;
14'd9396:data <=32'hFFAE003E;14'd9397:data <=32'hFFBF003A;14'd9398:data <=32'hFFC90031;
14'd9399:data <=32'hFFCB0024;14'd9400:data <=32'hFFC6001B;14'd9401:data <=32'hFFBB0016;
14'd9402:data <=32'hFFAE0017;14'd9403:data <=32'hFFA0001E;14'd9404:data <=32'hFF92002B;
14'd9405:data <=32'hFF87003E;14'd9406:data <=32'hFF7E0056;14'd9407:data <=32'hFF7A0074;
14'd9408:data <=32'hFFD2009E;14'd9409:data <=32'hFFDC00B3;14'd9410:data <=32'hFFE400B4;
14'd9411:data <=32'hFFA90096;14'd9412:data <=32'hFFBB00EE;14'd9413:data <=32'hFFEB0101;
14'd9414:data <=32'h00210105;14'd9415:data <=32'h005500FB;14'd9416:data <=32'h008300E4;
14'd9417:data <=32'h00A800C2;14'd9418:data <=32'h00C1009D;14'd9419:data <=32'h00D10076;
14'd9420:data <=32'h00D8004F;14'd9421:data <=32'h00DB002A;14'd9422:data <=32'h00D50006;
14'd9423:data <=32'h00CBFFE4;14'd9424:data <=32'h00BAFFC7;14'd9425:data <=32'h00A3FFAE;
14'd9426:data <=32'h0088FF9D;14'd9427:data <=32'h006DFF93;14'd9428:data <=32'h0053FF91;
14'd9429:data <=32'h003EFF96;14'd9430:data <=32'h002EFF9B;14'd9431:data <=32'h0022FFA2;
14'd9432:data <=32'h0018FFA6;14'd9433:data <=32'h000EFFA9;14'd9434:data <=32'h0003FFAE;
14'd9435:data <=32'hFFF7FFB4;14'd9436:data <=32'hFFECFFC0;14'd9437:data <=32'hFFE3FFD0;
14'd9438:data <=32'hFFE0FFE3;14'd9439:data <=32'hFFE6FFF6;14'd9440:data <=32'hFFF30005;
14'd9441:data <=32'h00060010;14'd9442:data <=32'h001B0012;14'd9443:data <=32'h0030000B;
14'd9444:data <=32'h0042FFFF;14'd9445:data <=32'h004FFFEC;14'd9446:data <=32'h0057FFD5;
14'd9447:data <=32'h0058FFBE;14'd9448:data <=32'h0054FFA5;14'd9449:data <=32'h0049FF8C;
14'd9450:data <=32'h0037FF74;14'd9451:data <=32'h001FFF62;14'd9452:data <=32'hFFFFFF54;
14'd9453:data <=32'hFFDCFF4F;14'd9454:data <=32'hFFB7FF56;14'd9455:data <=32'hFF95FF66;
14'd9456:data <=32'hFF79FF80;14'd9457:data <=32'hFF68FFA1;14'd9458:data <=32'hFF61FFC1;
14'd9459:data <=32'hFF67FFE0;14'd9460:data <=32'hFF73FFF8;14'd9461:data <=32'hFF820007;
14'd9462:data <=32'hFF92000E;14'd9463:data <=32'hFF9C000E;14'd9464:data <=32'hFFA1000C;
14'd9465:data <=32'hFFA3000A;14'd9466:data <=32'hFFA00009;14'd9467:data <=32'hFF9B000B;
14'd9468:data <=32'hFF95000F;14'd9469:data <=32'hFF8C0014;14'd9470:data <=32'hFF83001F;
14'd9471:data <=32'hFF7A002D;14'd9472:data <=32'hFF86FFEE;14'd9473:data <=32'hFF5F0006;
14'd9474:data <=32'hFF550029;14'd9475:data <=32'hFF9B0056;14'd9476:data <=32'hFF9B00A3;
14'd9477:data <=32'hFFBA00B0;14'd9478:data <=32'hFFDA00B6;14'd9479:data <=32'hFFF900B2;
14'd9480:data <=32'h001500A7;14'd9481:data <=32'h00270095;14'd9482:data <=32'h00320083;
14'd9483:data <=32'h00370075;14'd9484:data <=32'h0038006C;14'd9485:data <=32'h003B0067;
14'd9486:data <=32'h003F0064;14'd9487:data <=32'h00460060;14'd9488:data <=32'h0050005C;
14'd9489:data <=32'h00590055;14'd9490:data <=32'h0061004D;14'd9491:data <=32'h006A0044;
14'd9492:data <=32'h0072003A;14'd9493:data <=32'h007B002E;14'd9494:data <=32'h00830021;
14'd9495:data <=32'h008C000E;14'd9496:data <=32'h008EFFF6;14'd9497:data <=32'h008BFFDC;
14'd9498:data <=32'h007FFFC1;14'd9499:data <=32'h006BFFAA;14'd9500:data <=32'h004FFF9C;
14'd9501:data <=32'h002EFF98;14'd9502:data <=32'h0010FF9F;14'd9503:data <=32'hFFFAFFB1;
14'd9504:data <=32'hFFEAFFC7;14'd9505:data <=32'hFFE4FFE1;14'd9506:data <=32'hFFE9FFF9;
14'd9507:data <=32'hFFF4000C;14'd9508:data <=32'h0005001A;14'd9509:data <=32'h00180020;
14'd9510:data <=32'h002D0021;14'd9511:data <=32'h0043001C;14'd9512:data <=32'h00560012;
14'd9513:data <=32'h00670001;14'd9514:data <=32'h0074FFEA;14'd9515:data <=32'h007CFFCF;
14'd9516:data <=32'h0079FFB2;14'd9517:data <=32'h0070FF94;14'd9518:data <=32'h005DFF7B;
14'd9519:data <=32'h0045FF68;14'd9520:data <=32'h002AFF5D;14'd9521:data <=32'h000FFF5A;
14'd9522:data <=32'hFFF7FF5C;14'd9523:data <=32'hFFE3FF60;14'd9524:data <=32'hFFD4FF65;
14'd9525:data <=32'hFFC6FF69;14'd9526:data <=32'hFFB6FF6B;14'd9527:data <=32'hFFA3FF6D;
14'd9528:data <=32'hFF8CFF71;14'd9529:data <=32'hFF74FF7D;14'd9530:data <=32'hFF5DFF8E;
14'd9531:data <=32'hFF48FFA5;14'd9532:data <=32'hFF39FFC1;14'd9533:data <=32'hFF30FFE1;
14'd9534:data <=32'hFF2CFFFF;14'd9535:data <=32'hFF2E001F;14'd9536:data <=32'hFFDEFFAE;
14'd9537:data <=32'hFFAFFF9D;14'd9538:data <=32'hFF78FFAF;14'd9539:data <=32'hFF450050;
14'd9540:data <=32'hFF5000A8;14'd9541:data <=32'hFF7C00BD;14'd9542:data <=32'hFFAB00C5;
14'd9543:data <=32'hFFD800C0;14'd9544:data <=32'hFFFF00AC;14'd9545:data <=32'h00190090;
14'd9546:data <=32'h00270071;14'd9547:data <=32'h00270055;14'd9548:data <=32'h001E003F;
14'd9549:data <=32'h00110033;14'd9550:data <=32'h00040030;14'd9551:data <=32'hFFF70033;
14'd9552:data <=32'hFFF1003B;14'd9553:data <=32'hFFEE0044;14'd9554:data <=32'hFFEF0051;
14'd9555:data <=32'hFFF4005D;14'd9556:data <=32'hFFFD006A;14'd9557:data <=32'h000D0075;
14'd9558:data <=32'h0022007B;14'd9559:data <=32'h003B007B;14'd9560:data <=32'h00550073;
14'd9561:data <=32'h006D0062;14'd9562:data <=32'h007E0047;14'd9563:data <=32'h0085002B;
14'd9564:data <=32'h0082000D;14'd9565:data <=32'h0076FFF4;14'd9566:data <=32'h0065FFE2;
14'd9567:data <=32'h0051FFD9;14'd9568:data <=32'h003FFFD7;14'd9569:data <=32'h002FFFDA;
14'd9570:data <=32'h0024FFE0;14'd9571:data <=32'h001EFFE6;14'd9572:data <=32'h0019FFEE;
14'd9573:data <=32'h0016FFF4;14'd9574:data <=32'h0015FFFD;14'd9575:data <=32'h00150004;
14'd9576:data <=32'h0018000D;14'd9577:data <=32'h00200014;14'd9578:data <=32'h002B001A;
14'd9579:data <=32'h0037001C;14'd9580:data <=32'h0046001A;14'd9581:data <=32'h00540014;
14'd9582:data <=32'h0060000A;14'd9583:data <=32'h006BFFFF;14'd9584:data <=32'h0073FFF1;
14'd9585:data <=32'h007CFFE4;14'd9586:data <=32'h0084FFD3;14'd9587:data <=32'h008CFFBE;
14'd9588:data <=32'h0092FFA4;14'd9589:data <=32'h0093FF83;14'd9590:data <=32'h008AFF5D;
14'd9591:data <=32'h0075FF35;14'd9592:data <=32'h0053FF11;14'd9593:data <=32'h0026FEF5;
14'd9594:data <=32'hFFF0FEE5;14'd9595:data <=32'hFFB6FEE5;14'd9596:data <=32'hFF7EFEF3;
14'd9597:data <=32'hFF4AFF0F;14'd9598:data <=32'hFF1FFF35;14'd9599:data <=32'hFEFDFF63;
14'd9600:data <=32'hFFD2FFAB;14'd9601:data <=32'hFFB7FF95;14'd9602:data <=32'hFF87FF7F;
14'd9603:data <=32'hFEF9FF94;14'd9604:data <=32'hFEE30005;14'd9605:data <=32'hFEF9003A;
14'd9606:data <=32'hFF1B0065;14'd9607:data <=32'hFF440085;14'd9608:data <=32'hFF700092;
14'd9609:data <=32'hFF990093;14'd9610:data <=32'hFFBB008A;14'd9611:data <=32'hFFD1007B;
14'd9612:data <=32'hFFDF006B;14'd9613:data <=32'hFFE6005E;14'd9614:data <=32'hFFE90055;
14'd9615:data <=32'hFFEA004F;14'd9616:data <=32'hFFEC004C;14'd9617:data <=32'hFFEE0049;
14'd9618:data <=32'hFFEF0046;14'd9619:data <=32'hFFEF0045;14'd9620:data <=32'hFFEF0047;
14'd9621:data <=32'hFFF0004B;14'd9622:data <=32'hFFF30050;14'd9623:data <=32'hFFFA0055;
14'd9624:data <=32'h00060058;14'd9625:data <=32'h00120057;14'd9626:data <=32'h001D0052;
14'd9627:data <=32'h0025004A;14'd9628:data <=32'h0029003F;14'd9629:data <=32'h00290037;
14'd9630:data <=32'h00250031;14'd9631:data <=32'h00220031;14'd9632:data <=32'h00210033;
14'd9633:data <=32'h00260037;14'd9634:data <=32'h002C0039;14'd9635:data <=32'h00360037;
14'd9636:data <=32'h00400030;14'd9637:data <=32'h00470026;14'd9638:data <=32'h0049001A;
14'd9639:data <=32'h0047000F;14'd9640:data <=32'h00400005;14'd9641:data <=32'h00370000;
14'd9642:data <=32'h002EFFFF;14'd9643:data <=32'h00260002;14'd9644:data <=32'h00210007;
14'd9645:data <=32'h001D000F;14'd9646:data <=32'h001D0019;14'd9647:data <=32'h00210023;
14'd9648:data <=32'h002A002F;14'd9649:data <=32'h0038003A;14'd9650:data <=32'h004D0043;
14'd9651:data <=32'h00690046;14'd9652:data <=32'h008B003E;14'd9653:data <=32'h00AC002B;
14'd9654:data <=32'h00CB000A;14'd9655:data <=32'h00E0FFDC;14'd9656:data <=32'h00E7FFA7;
14'd9657:data <=32'h00DDFF6F;14'd9658:data <=32'h00C4FF3C;14'd9659:data <=32'h009CFF10;
14'd9660:data <=32'h006CFEF1;14'd9661:data <=32'h0036FEDE;14'd9662:data <=32'hFFFFFED8;
14'd9663:data <=32'hFFC9FEDE;14'd9664:data <=32'hFFFDFF31;14'd9665:data <=32'hFFD7FF18;
14'd9666:data <=32'hFFB8FF04;14'd9667:data <=32'hFFB5FEF0;14'd9668:data <=32'hFF78FF3F;
14'd9669:data <=32'hFF62FF5D;14'd9670:data <=32'hFF54FF7E;14'd9671:data <=32'hFF4EFF9D;
14'd9672:data <=32'hFF4EFFB8;14'd9673:data <=32'hFF52FFCC;14'd9674:data <=32'hFF53FFDD;
14'd9675:data <=32'hFF53FFED;14'd9676:data <=32'hFF52FFFE;14'd9677:data <=32'hFF500013;
14'd9678:data <=32'hFF53002A;14'd9679:data <=32'hFF5C0046;14'd9680:data <=32'hFF6B005F;
14'd9681:data <=32'hFF820073;14'd9682:data <=32'hFF9D0080;14'd9683:data <=32'hFFB90086;
14'd9684:data <=32'hFFD20084;14'd9685:data <=32'hFFEA007E;14'd9686:data <=32'hFFFE0075;
14'd9687:data <=32'h000E0068;14'd9688:data <=32'h001C0059;14'd9689:data <=32'h00250047;
14'd9690:data <=32'h00290033;14'd9691:data <=32'h0026001F;14'd9692:data <=32'h001B000D;
14'd9693:data <=32'h000B0000;14'd9694:data <=32'hFFF7FFFC;14'd9695:data <=32'hFFE10001;
14'd9696:data <=32'hFFD20010;14'd9697:data <=32'hFFC90025;14'd9698:data <=32'hFFC9003B;
14'd9699:data <=32'hFFD3004F;14'd9700:data <=32'hFFE3005E;14'd9701:data <=32'hFFF60065;
14'd9702:data <=32'h00080066;14'd9703:data <=32'h00190062;14'd9704:data <=32'h0025005A;
14'd9705:data <=32'h002E0051;14'd9706:data <=32'h00340048;14'd9707:data <=32'h0037003F;
14'd9708:data <=32'h00380039;14'd9709:data <=32'h00370034;14'd9710:data <=32'h00360030;
14'd9711:data <=32'h0034002F;14'd9712:data <=32'h00320031;14'd9713:data <=32'h00330036;
14'd9714:data <=32'h0037003F;14'd9715:data <=32'h00430049;14'd9716:data <=32'h0055004F;
14'd9717:data <=32'h006C004F;14'd9718:data <=32'h00870046;14'd9719:data <=32'h00A10033;
14'd9720:data <=32'h00B40017;14'd9721:data <=32'h00BFFFF5;14'd9722:data <=32'h00C0FFD2;
14'd9723:data <=32'h00B7FFB0;14'd9724:data <=32'h00A8FF93;14'd9725:data <=32'h0094FF7C;
14'd9726:data <=32'h007FFF6A;14'd9727:data <=32'h006AFF5C;14'd9728:data <=32'h00CBFF42;
14'd9729:data <=32'h00B0FF06;14'd9730:data <=32'h0088FEE9;14'd9731:data <=32'h0068FF55;
14'd9732:data <=32'h003FFF80;14'd9733:data <=32'h0038FF77;14'd9734:data <=32'h002FFF6F;
14'd9735:data <=32'h0024FF64;14'd9736:data <=32'h0017FF57;14'd9737:data <=32'h0005FF48;
14'd9738:data <=32'hFFEDFF3B;14'd9739:data <=32'hFFCCFF31;14'd9740:data <=32'hFFA3FF31;
14'd9741:data <=32'hFF77FF3D;14'd9742:data <=32'hFF4EFF57;14'd9743:data <=32'hFF2DFF7D;
14'd9744:data <=32'hFF18FFAC;14'd9745:data <=32'hFF11FFDE;14'd9746:data <=32'hFF18000E;
14'd9747:data <=32'hFF2A0039;14'd9748:data <=32'hFF44005D;14'd9749:data <=32'hFF650077;
14'd9750:data <=32'hFF880088;14'd9751:data <=32'hFFAE0091;14'd9752:data <=32'hFFD10090;
14'd9753:data <=32'hFFF50087;14'd9754:data <=32'h00140074;14'd9755:data <=32'h00280058;
14'd9756:data <=32'h0034003A;14'd9757:data <=32'h00340019;14'd9758:data <=32'h0028FFFE;
14'd9759:data <=32'h0015FFE9;14'd9760:data <=32'hFFFDFFDF;14'd9761:data <=32'hFFE4FFDF;
14'd9762:data <=32'hFFCFFFE7;14'd9763:data <=32'hFFC0FFF3;14'd9764:data <=32'hFFB70003;
14'd9765:data <=32'hFFB30013;14'd9766:data <=32'hFFB10020;14'd9767:data <=32'hFFB1002D;
14'd9768:data <=32'hFFB1003A;14'd9769:data <=32'hFFB30046;14'd9770:data <=32'hFFB70056;
14'd9771:data <=32'hFFBE0066;14'd9772:data <=32'hFFC90076;14'd9773:data <=32'hFFD80084;
14'd9774:data <=32'hFFEA008F;14'd9775:data <=32'hFFFF0095;14'd9776:data <=32'h0014009A;
14'd9777:data <=32'h00290099;14'd9778:data <=32'h003F0097;14'd9779:data <=32'h00550093;
14'd9780:data <=32'h006C008B;14'd9781:data <=32'h0085007E;14'd9782:data <=32'h009C0069;
14'd9783:data <=32'h00AF004F;14'd9784:data <=32'h00BB002E;14'd9785:data <=32'h00BD000B;
14'd9786:data <=32'h00B4FFE8;14'd9787:data <=32'h00A2FFCE;14'd9788:data <=32'h008AFFBB;
14'd9789:data <=32'h0073FFB3;14'd9790:data <=32'h005EFFB3;14'd9791:data <=32'h0050FFB9;
14'd9792:data <=32'h00F1000F;14'd9793:data <=32'h0109FFD8;14'd9794:data <=32'h00F9FF9E;
14'd9795:data <=32'h0062FFB0;14'd9796:data <=32'h0048FFE7;14'd9797:data <=32'h0053FFE7;
14'd9798:data <=32'h0062FFE3;14'd9799:data <=32'h0070FFD6;14'd9800:data <=32'h007DFFC4;
14'd9801:data <=32'h0084FFA8;14'd9802:data <=32'h0084FF85;14'd9803:data <=32'h0077FF62;
14'd9804:data <=32'h005CFF3F;14'd9805:data <=32'h0035FF24;14'd9806:data <=32'h0007FF19;
14'd9807:data <=32'hFFD6FF1B;14'd9808:data <=32'hFFA8FF2A;14'd9809:data <=32'hFF83FF45;
14'd9810:data <=32'hFF67FF65;14'd9811:data <=32'hFF56FF89;14'd9812:data <=32'hFF4DFFAD;
14'd9813:data <=32'hFF4CFFD1;14'd9814:data <=32'hFF51FFF2;14'd9815:data <=32'hFF5C0010;
14'd9816:data <=32'hFF6D002A;14'd9817:data <=32'hFF830040;14'd9818:data <=32'hFF9E004D;
14'd9819:data <=32'hFFBA0053;14'd9820:data <=32'hFFD50050;14'd9821:data <=32'hFFEA0046;
14'd9822:data <=32'hFFFA0036;14'd9823:data <=32'h00020026;14'd9824:data <=32'h00050017;
14'd9825:data <=32'h0004000B;14'd9826:data <=32'h00020001;14'd9827:data <=32'hFFFFFFF8;
14'd9828:data <=32'hFFFBFFEE;14'd9829:data <=32'hFFF5FFE3;14'd9830:data <=32'hFFEBFFD9;
14'd9831:data <=32'hFFDCFFCE;14'd9832:data <=32'hFFC8FFC8;14'd9833:data <=32'hFFAEFFC8;
14'd9834:data <=32'hFF94FFD1;14'd9835:data <=32'hFF78FFE4;14'd9836:data <=32'hFF64FFFF;
14'd9837:data <=32'hFF570022;14'd9838:data <=32'hFF530048;14'd9839:data <=32'hFF59006E;
14'd9840:data <=32'hFF680093;14'd9841:data <=32'hFF7F00B5;14'd9842:data <=32'hFFA000D2;
14'd9843:data <=32'hFFC500E9;14'd9844:data <=32'hFFF100F8;14'd9845:data <=32'h002100FC;
14'd9846:data <=32'h005400F3;14'd9847:data <=32'h008300DE;14'd9848:data <=32'h00AB00BC;
14'd9849:data <=32'h00C70090;14'd9850:data <=32'h00D5005F;14'd9851:data <=32'h00D40030;
14'd9852:data <=32'h00C40008;14'd9853:data <=32'h00ADFFEA;14'd9854:data <=32'h0093FFD8;
14'd9855:data <=32'h007AFFD1;14'd9856:data <=32'h0078004B;14'd9857:data <=32'h00950042;
14'd9858:data <=32'h00B0001E;14'd9859:data <=32'h009CFFC8;14'd9860:data <=32'h0075FFF4;
14'd9861:data <=32'h0074FFF0;14'd9862:data <=32'h0074FFEB;14'd9863:data <=32'h0076FFE5;
14'd9864:data <=32'h007BFFDD;14'd9865:data <=32'h007FFFD0;14'd9866:data <=32'h0083FFBE;
14'd9867:data <=32'h0080FFA7;14'd9868:data <=32'h0076FF90;14'd9869:data <=32'h0062FF79;
14'd9870:data <=32'h0049FF6A;14'd9871:data <=32'h002CFF64;14'd9872:data <=32'h0010FF67;
14'd9873:data <=32'hFFF9FF70;14'd9874:data <=32'hFFE9FF7D;14'd9875:data <=32'hFFDEFF8A;
14'd9876:data <=32'hFFD7FF95;14'd9877:data <=32'hFFD2FF9D;14'd9878:data <=32'hFFCCFFA5;
14'd9879:data <=32'hFFC5FFAC;14'd9880:data <=32'hFFBFFFB3;14'd9881:data <=32'hFFBAFFBD;
14'd9882:data <=32'hFFB6FFC8;14'd9883:data <=32'hFFB5FFD2;14'd9884:data <=32'hFFB5FFDC;
14'd9885:data <=32'hFFB7FFE5;14'd9886:data <=32'hFFB8FFEC;14'd9887:data <=32'hFFB9FFF3;
14'd9888:data <=32'hFFBBFFFC;14'd9889:data <=32'hFFC00006;14'd9890:data <=32'hFFC80010;
14'd9891:data <=32'hFFD50018;14'd9892:data <=32'hFFE6001A;14'd9893:data <=32'hFFF80014;
14'd9894:data <=32'h00080007;14'd9895:data <=32'h0012FFF2;14'd9896:data <=32'h0012FFD8;
14'd9897:data <=32'h0007FFBF;14'd9898:data <=32'hFFF2FFA9;14'd9899:data <=32'hFFD5FF9B;
14'd9900:data <=32'hFFB3FF98;14'd9901:data <=32'hFF91FF9F;14'd9902:data <=32'hFF71FFB1;
14'd9903:data <=32'hFF56FFCA;14'd9904:data <=32'hFF41FFEA;14'd9905:data <=32'hFF34000F;
14'd9906:data <=32'hFF2F0037;14'd9907:data <=32'hFF340062;14'd9908:data <=32'hFF42008B;
14'd9909:data <=32'hFF5B00B2;14'd9910:data <=32'hFF7E00D3;14'd9911:data <=32'hFFAA00E9;
14'd9912:data <=32'hFFD800F2;14'd9913:data <=32'h000400EE;14'd9914:data <=32'h002C00E0;
14'd9915:data <=32'h004A00CB;14'd9916:data <=32'h006000B3;14'd9917:data <=32'h006D009E;
14'd9918:data <=32'h0076008A;14'd9919:data <=32'h007C007C;14'd9920:data <=32'h00710041;
14'd9921:data <=32'h0076003C;14'd9922:data <=32'h00850041;14'd9923:data <=32'h00B9007F;
14'd9924:data <=32'h00AF0096;14'd9925:data <=32'h00C60079;14'd9926:data <=32'h00D60058;
14'd9927:data <=32'h00DF0033;14'd9928:data <=32'h00E10010;14'd9929:data <=32'h00DDFFEC;
14'd9930:data <=32'h00D5FFC7;14'd9931:data <=32'h00C3FFA5;14'd9932:data <=32'h00AAFF86;
14'd9933:data <=32'h0089FF6E;14'd9934:data <=32'h0062FF61;14'd9935:data <=32'h0039FF60;
14'd9936:data <=32'h0014FF6A;14'd9937:data <=32'hFFF8FF7F;14'd9938:data <=32'hFFE8FF9B;
14'd9939:data <=32'hFFE2FFB5;14'd9940:data <=32'hFFE7FFCC;14'd9941:data <=32'hFFF1FFDB;
14'd9942:data <=32'hFFFFFFE3;14'd9943:data <=32'h000BFFE3;14'd9944:data <=32'h0014FFDF;
14'd9945:data <=32'h001BFFD7;14'd9946:data <=32'h001DFFD0;14'd9947:data <=32'h001DFFC6;
14'd9948:data <=32'h001AFFBC;14'd9949:data <=32'h0013FFB2;14'd9950:data <=32'h0008FFAA;
14'd9951:data <=32'hFFFAFFA6;14'd9952:data <=32'hFFEAFFA5;14'd9953:data <=32'hFFDAFFAC;
14'd9954:data <=32'hFFCDFFB7;14'd9955:data <=32'hFFC6FFC8;14'd9956:data <=32'hFFC6FFD8;
14'd9957:data <=32'hFFCEFFE6;14'd9958:data <=32'hFFD9FFEE;14'd9959:data <=32'hFFE7FFEF;
14'd9960:data <=32'hFFF3FFE7;14'd9961:data <=32'hFFF9FFDB;14'd9962:data <=32'hFFF9FFCD;
14'd9963:data <=32'hFFF1FFBF;14'd9964:data <=32'hFFE4FFB5;14'd9965:data <=32'hFFD6FFAF;
14'd9966:data <=32'hFFC5FFAE;14'd9967:data <=32'hFFB5FFB0;14'd9968:data <=32'hFFA5FFB5;
14'd9969:data <=32'hFF97FFBD;14'd9970:data <=32'hFF88FFC7;14'd9971:data <=32'hFF7AFFD4;
14'd9972:data <=32'hFF6DFFE4;14'd9973:data <=32'hFF63FFF9;14'd9974:data <=32'hFF5F000F;
14'd9975:data <=32'hFF5F0026;14'd9976:data <=32'hFF63003B;14'd9977:data <=32'hFF6B004F;
14'd9978:data <=32'hFF71005F;14'd9979:data <=32'hFF77006E;14'd9980:data <=32'hFF7D007E;
14'd9981:data <=32'hFF830093;14'd9982:data <=32'hFF8B00AB;14'd9983:data <=32'hFF9D00C8;
14'd9984:data <=32'h003700A1;14'd9985:data <=32'h0044009E;14'd9986:data <=32'h003E009D;
14'd9987:data <=32'hFFE100F3;14'd9988:data <=32'hFFF30130;14'd9989:data <=32'h002F0130;
14'd9990:data <=32'h00690123;14'd9991:data <=32'h009D0107;14'd9992:data <=32'h00CA00E2;
14'd9993:data <=32'h00EE00B5;14'd9994:data <=32'h01070080;14'd9995:data <=32'h01140047;
14'd9996:data <=32'h0112000C;14'd9997:data <=32'h0101FFD4;14'd9998:data <=32'h00E1FFA5;
14'd9999:data <=32'h00B6FF82;14'd10000:data <=32'h0086FF70;14'd10001:data <=32'h0058FF6D;
14'd10002:data <=32'h0030FF78;14'd10003:data <=32'h0012FF8B;14'd10004:data <=32'hFFFFFFA4;
14'd10005:data <=32'hFFF7FFBA;14'd10006:data <=32'hFFF5FFCE;14'd10007:data <=32'hFFF8FFDE;
14'd10008:data <=32'hFFFEFFE9;14'd10009:data <=32'h0005FFF3;14'd10010:data <=32'h000EFFF9;
14'd10011:data <=32'h0018FFFC;14'd10012:data <=32'h0023FFFC;14'd10013:data <=32'h002EFFF6;
14'd10014:data <=32'h0037FFEE;14'd10015:data <=32'h003BFFE3;14'd10016:data <=32'h003BFFD7;
14'd10017:data <=32'h0037FFCB;14'd10018:data <=32'h0031FFC3;14'd10019:data <=32'h0029FFBD;
14'd10020:data <=32'h0024FFBA;14'd10021:data <=32'h0020FFB8;14'd10022:data <=32'h001DFFB4;
14'd10023:data <=32'h001BFFAD;14'd10024:data <=32'h0017FFA4;14'd10025:data <=32'h000EFF9B;
14'd10026:data <=32'h0000FF91;14'd10027:data <=32'hFFEFFF8D;14'd10028:data <=32'hFFDAFF8E;
14'd10029:data <=32'hFFC7FF95;14'd10030:data <=32'hFFB9FFA2;14'd10031:data <=32'hFFAFFFB3;
14'd10032:data <=32'hFFACFFC1;14'd10033:data <=32'hFFAEFFCF;14'd10034:data <=32'hFFB3FFD8;
14'd10035:data <=32'hFFB8FFDD;14'd10036:data <=32'hFFBCFFDF;14'd10037:data <=32'hFFBFFFDD;
14'd10038:data <=32'hFFBFFFDA;14'd10039:data <=32'hFFBDFFD6;14'd10040:data <=32'hFFB9FFCF;
14'd10041:data <=32'hFFB0FFC9;14'd10042:data <=32'hFFA1FFC2;14'd10043:data <=32'hFF8BFFC0;
14'd10044:data <=32'hFF70FFC3;14'd10045:data <=32'hFF4FFFD1;14'd10046:data <=32'hFF31FFED;
14'd10047:data <=32'hFF180016;14'd10048:data <=32'hFF7A0068;14'd10049:data <=32'hFF770083;
14'd10050:data <=32'hFF7B0088;14'd10051:data <=32'hFF41005E;14'd10052:data <=32'hFF3200B8;
14'd10053:data <=32'hFF5700DE;14'd10054:data <=32'hFF8300FA;14'd10055:data <=32'hFFB4010A;
14'd10056:data <=32'hFFE50111;14'd10057:data <=32'h0016010E;14'd10058:data <=32'h00470101;
14'd10059:data <=32'h007100E9;14'd10060:data <=32'h009600C8;14'd10061:data <=32'h00B0009F;
14'd10062:data <=32'h00BE0073;14'd10063:data <=32'h00BF004A;14'd10064:data <=32'h00B50025;
14'd10065:data <=32'h00A50009;14'd10066:data <=32'h0092FFF5;14'd10067:data <=32'h0081FFE9;
14'd10068:data <=32'h0073FFE1;14'd10069:data <=32'h0068FFDA;14'd10070:data <=32'h005EFFD3;
14'd10071:data <=32'h0052FFCC;14'd10072:data <=32'h0043FFC5;14'd10073:data <=32'h0034FFC3;
14'd10074:data <=32'h0023FFC5;14'd10075:data <=32'h0015FFCC;14'd10076:data <=32'h0009FFD7;
14'd10077:data <=32'h0004FFE5;14'd10078:data <=32'h0002FFF3;14'd10079:data <=32'h0006FFFF;
14'd10080:data <=32'h000D0009;14'd10081:data <=32'h00160011;14'd10082:data <=32'h00210017;
14'd10083:data <=32'h002F001B;14'd10084:data <=32'h003F001B;14'd10085:data <=32'h00500015;
14'd10086:data <=32'h0063000A;14'd10087:data <=32'h0074FFF7;14'd10088:data <=32'h007FFFDD;
14'd10089:data <=32'h0081FFBD;14'd10090:data <=32'h0079FF9E;14'd10091:data <=32'h0067FF80;
14'd10092:data <=32'h004CFF6A;14'd10093:data <=32'h002CFF5D;14'd10094:data <=32'h000AFF5C;
14'd10095:data <=32'hFFECFF63;14'd10096:data <=32'hFFD5FF72;14'd10097:data <=32'hFFC5FF84;
14'd10098:data <=32'hFFBBFF97;14'd10099:data <=32'hFFB9FFA7;14'd10100:data <=32'hFFB9FFB5;
14'd10101:data <=32'hFFBBFFBF;14'd10102:data <=32'hFFC0FFC6;14'd10103:data <=32'hFFC5FFCA;
14'd10104:data <=32'hFFCBFFC9;14'd10105:data <=32'hFFD0FFC3;14'd10106:data <=32'hFFCEFFB9;
14'd10107:data <=32'hFFC7FFAB;14'd10108:data <=32'hFFB7FF9E;14'd10109:data <=32'hFF9EFF97;
14'd10110:data <=32'hFF7FFF99;14'd10111:data <=32'hFF5DFFA7;14'd10112:data <=32'hFF82FF94;
14'd10113:data <=32'hFF51FF9F;14'd10114:data <=32'hFF3AFFBB;14'd10115:data <=32'hFF6AFFF1;
14'd10116:data <=32'hFF470038;14'd10117:data <=32'hFF570051;14'd10118:data <=32'hFF690065;
14'd10119:data <=32'hFF7D0072;14'd10120:data <=32'hFF8F007C;14'd10121:data <=32'hFFA00085;
14'd10122:data <=32'hFFB2008C;14'd10123:data <=32'hFFC40091;14'd10124:data <=32'hFFD60092;
14'd10125:data <=32'hFFE80091;14'd10126:data <=32'hFFF6008C;14'd10127:data <=32'h00020088;
14'd10128:data <=32'h000B0085;14'd10129:data <=32'h00140084;14'd10130:data <=32'h001F0085;
14'd10131:data <=32'h002E0087;14'd10132:data <=32'h00420086;14'd10133:data <=32'h0059007E;
14'd10134:data <=32'h0071006F;14'd10135:data <=32'h00840057;14'd10136:data <=32'h008F0039;
14'd10137:data <=32'h00900019;14'd10138:data <=32'h0087FFFA;14'd10139:data <=32'h0076FFE2;
14'd10140:data <=32'h0060FFD1;14'd10141:data <=32'h0047FFC8;14'd10142:data <=32'h0030FFC7;
14'd10143:data <=32'h001AFFCB;14'd10144:data <=32'h0007FFD5;14'd10145:data <=32'hFFF8FFE6;
14'd10146:data <=32'hFFF0FFF8;14'd10147:data <=32'hFFED000E;14'd10148:data <=32'hFFF20025;
14'd10149:data <=32'h0000003B;14'd10150:data <=32'h0016004A;14'd10151:data <=32'h00320053;
14'd10152:data <=32'h00510051;14'd10153:data <=32'h006E0043;14'd10154:data <=32'h0085002C;
14'd10155:data <=32'h0095000F;14'd10156:data <=32'h009AFFF0;14'd10157:data <=32'h0096FFD3;
14'd10158:data <=32'h008CFFBA;14'd10159:data <=32'h007EFFA8;14'd10160:data <=32'h0070FF99;
14'd10161:data <=32'h0063FF8D;14'd10162:data <=32'h0055FF83;14'd10163:data <=32'h0048FF78;
14'd10164:data <=32'h003AFF6F;14'd10165:data <=32'h002AFF66;14'd10166:data <=32'h0018FF60;
14'd10167:data <=32'h0005FF5C;14'd10168:data <=32'hFFF2FF5A;14'd10169:data <=32'hFFDFFF5B;
14'd10170:data <=32'hFFCCFF5D;14'd10171:data <=32'hFFBAFF60;14'd10172:data <=32'hFFA5FF64;
14'd10173:data <=32'hFF8CFF6B;14'd10174:data <=32'hFF74FF77;14'd10175:data <=32'hFF5BFF8B;
14'd10176:data <=32'h001AFF71;14'd10177:data <=32'hFFEEFF4D;14'd10178:data <=32'hFFB3FF4A;
14'd10179:data <=32'hFF52FFD2;14'd10180:data <=32'hFF380022;14'd10181:data <=32'hFF54003E;
14'd10182:data <=32'hFF73004E;14'd10183:data <=32'hFF920055;14'd10184:data <=32'hFFAA0051;
14'd10185:data <=32'hFFBC0048;14'd10186:data <=32'hFFC7003F;14'd10187:data <=32'hFFCE0035;
14'd10188:data <=32'hFFCF002C;14'd10189:data <=32'hFFCD0024;14'd10190:data <=32'hFFC6001E;
14'd10191:data <=32'hFFBB001F;14'd10192:data <=32'hFFB00023;14'd10193:data <=32'hFFA30030;
14'd10194:data <=32'hFF9B0045;14'd10195:data <=32'hFF9C005F;14'd10196:data <=32'hFFA7007B;
14'd10197:data <=32'hFFBD0092;14'd10198:data <=32'hFFDD00A3;14'd10199:data <=32'hFFFF00A8;
14'd10200:data <=32'h002300A0;14'd10201:data <=32'h00400090;14'd10202:data <=32'h00560079;
14'd10203:data <=32'h00630060;14'd10204:data <=32'h00670045;14'd10205:data <=32'h0066002D;
14'd10206:data <=32'h00600019;14'd10207:data <=32'h00560008;14'd10208:data <=32'h0049FFFA;
14'd10209:data <=32'h003AFFF1;14'd10210:data <=32'h002AFFEC;14'd10211:data <=32'h0016FFED;
14'd10212:data <=32'h0007FFF5;14'd10213:data <=32'hFFFB0002;14'd10214:data <=32'hFFF50013;
14'd10215:data <=32'hFFF60024;14'd10216:data <=32'hFFFE0035;14'd10217:data <=32'h00090041;
14'd10218:data <=32'h00180048;14'd10219:data <=32'h0027004A;14'd10220:data <=32'h0035004B;
14'd10221:data <=32'h0041004A;14'd10222:data <=32'h004D0049;14'd10223:data <=32'h005B0049;
14'd10224:data <=32'h006E0048;14'd10225:data <=32'h00850040;14'd10226:data <=32'h009D0033;
14'd10227:data <=32'h00B5001F;14'd10228:data <=32'h00C9FFFF;14'd10229:data <=32'h00D6FFD9;
14'd10230:data <=32'h00D9FFAE;14'd10231:data <=32'h00D1FF83;14'd10232:data <=32'h00BFFF58;
14'd10233:data <=32'h00A3FF32;14'd10234:data <=32'h0080FF12;14'd10235:data <=32'h0057FEF9;
14'd10236:data <=32'h0028FEE7;14'd10237:data <=32'hFFF2FEDF;14'd10238:data <=32'hFFBBFEE4;
14'd10239:data <=32'hFF85FEF7;14'd10240:data <=32'h002EFF97;14'd10241:data <=32'h001EFF70;
14'd10242:data <=32'hFFF8FF47;14'd10243:data <=32'hFF61FF2E;14'd10244:data <=32'hFF25FF89;
14'd10245:data <=32'hFF29FFBA;14'd10246:data <=32'hFF37FFE4;14'd10247:data <=32'hFF4E0003;
14'd10248:data <=32'hFF660017;14'd10249:data <=32'hFF7D0022;14'd10250:data <=32'hFF910028;
14'd10251:data <=32'hFFA3002A;14'd10252:data <=32'hFFB10026;14'd10253:data <=32'hFFBC0022;
14'd10254:data <=32'hFFC3001A;14'd10255:data <=32'hFFC40011;14'd10256:data <=32'hFFC1000B;
14'd10257:data <=32'hFFB70008;14'd10258:data <=32'hFFAC000C;14'd10259:data <=32'hFFA10017;
14'd10260:data <=32'hFF9D0028;14'd10261:data <=32'hFF9F003C;14'd10262:data <=32'hFFAA004D;
14'd10263:data <=32'hFFB9005A;14'd10264:data <=32'hFFCB0061;14'd10265:data <=32'hFFDC0061;
14'd10266:data <=32'hFFEA005D;14'd10267:data <=32'hFFF20057;14'd10268:data <=32'hFFF90052;
14'd10269:data <=32'hFFFD004F;14'd10270:data <=32'h0001004E;14'd10271:data <=32'h0008004C;
14'd10272:data <=32'h000F004B;14'd10273:data <=32'h00160046;14'd10274:data <=32'h001C0040;
14'd10275:data <=32'h001E0038;14'd10276:data <=32'h00200032;14'd10277:data <=32'h001F002B;
14'd10278:data <=32'h001E0025;14'd10279:data <=32'h001A0022;14'd10280:data <=32'h0018001F;
14'd10281:data <=32'h0015001D;14'd10282:data <=32'h0010001A;14'd10283:data <=32'h0009001A;
14'd10284:data <=32'h0000001D;14'd10285:data <=32'hFFF60025;14'd10286:data <=32'hFFED0034;
14'd10287:data <=32'hFFE90049;14'd10288:data <=32'hFFEF0064;14'd10289:data <=32'h0000007E;
14'd10290:data <=32'h001D0095;14'd10291:data <=32'h004400A3;14'd10292:data <=32'h007000A4;
14'd10293:data <=32'h009F0098;14'd10294:data <=32'h00C9007E;14'd10295:data <=32'h00EC0059;
14'd10296:data <=32'h0106002B;14'd10297:data <=32'h0114FFF9;14'd10298:data <=32'h0118FFC2;
14'd10299:data <=32'h010EFF8B;14'd10300:data <=32'h00F9FF56;14'd10301:data <=32'h00D8FF25;
14'd10302:data <=32'h00A9FEFC;14'd10303:data <=32'h0071FEE0;14'd10304:data <=32'h006EFF59;
14'd10305:data <=32'h005AFF34;14'd10306:data <=32'h004BFF14;14'd10307:data <=32'h0048FEEE;
14'd10308:data <=32'hFFF3FF1F;14'd10309:data <=32'hFFD8FF31;14'd10310:data <=32'hFFC5FF42;
14'd10311:data <=32'hFFB6FF52;14'd10312:data <=32'hFFA9FF60;14'd10313:data <=32'hFF9AFF6C;
14'd10314:data <=32'hFF8BFF7A;14'd10315:data <=32'hFF7DFF8C;14'd10316:data <=32'hFF72FFA0;
14'd10317:data <=32'hFF6AFFB6;14'd10318:data <=32'hFF68FFCD;14'd10319:data <=32'hFF69FFE1;
14'd10320:data <=32'hFF6DFFF4;14'd10321:data <=32'hFF720006;14'd10322:data <=32'hFF780017;
14'd10323:data <=32'hFF810029;14'd10324:data <=32'hFF8E0039;14'd10325:data <=32'hFFA00047;
14'd10326:data <=32'hFFB50051;14'd10327:data <=32'hFFCD0053;14'd10328:data <=32'hFFE3004C;
14'd10329:data <=32'hFFF5003E;14'd10330:data <=32'hFFFF002B;14'd10331:data <=32'h00000018;
14'd10332:data <=32'hFFF60008;14'd10333:data <=32'hFFE9FFFF;14'd10334:data <=32'hFFD9FFFD;
14'd10335:data <=32'hFFCB0003;14'd10336:data <=32'hFFC2000D;14'd10337:data <=32'hFFBD001A;
14'd10338:data <=32'hFFBC0028;14'd10339:data <=32'hFFBF0033;14'd10340:data <=32'hFFC5003E;
14'd10341:data <=32'hFFCD0048;14'd10342:data <=32'hFFD8004F;14'd10343:data <=32'hFFE30053;
14'd10344:data <=32'hFFF00054;14'd10345:data <=32'hFFFC0052;14'd10346:data <=32'h0006004A;
14'd10347:data <=32'h000C0040;14'd10348:data <=32'h000B0036;14'd10349:data <=32'h0005002D;
14'd10350:data <=32'hFFFA002A;14'd10351:data <=32'hFFEC002F;14'd10352:data <=32'hFFE1003D;
14'd10353:data <=32'hFFDD0052;14'd10354:data <=32'hFFE1006A;14'd10355:data <=32'hFFF10082;
14'd10356:data <=32'h00090095;14'd10357:data <=32'h002700A0;14'd10358:data <=32'h004800A1;
14'd10359:data <=32'h0069009B;14'd10360:data <=32'h0087008D;14'd10361:data <=32'h00A20079;
14'd10362:data <=32'h00B90061;14'd10363:data <=32'h00CB0045;14'd10364:data <=32'h00D90024;
14'd10365:data <=32'h00DF0000;14'd10366:data <=32'h00DFFFDA;14'd10367:data <=32'h00D6FFB6;
14'd10368:data <=32'h0112FFBA;14'd10369:data <=32'h0111FF7B;14'd10370:data <=32'h00FAFF58;
14'd10371:data <=32'h00C8FFAC;14'd10372:data <=32'h0094FFC3;14'd10373:data <=32'h0097FFB6;
14'd10374:data <=32'h009AFFA2;14'd10375:data <=32'h009AFF8A;14'd10376:data <=32'h0093FF6A;
14'd10377:data <=32'h0080FF4A;14'd10378:data <=32'h0065FF2C;14'd10379:data <=32'h003EFF17;
14'd10380:data <=32'h0011FF0B;14'd10381:data <=32'hFFE3FF0B;14'd10382:data <=32'hFFB7FF17;
14'd10383:data <=32'hFF90FF2C;14'd10384:data <=32'hFF6EFF48;14'd10385:data <=32'hFF53FF69;
14'd10386:data <=32'hFF40FF91;14'd10387:data <=32'hFF36FFBB;14'd10388:data <=32'hFF37FFE8;
14'd10389:data <=32'hFF420012;14'd10390:data <=32'hFF5A0038;14'd10391:data <=32'hFF7C0054;
14'd10392:data <=32'hFFA30062;14'd10393:data <=32'hFFCB0063;14'd10394:data <=32'hFFED0056;
14'd10395:data <=32'h00060041;14'd10396:data <=32'h00140026;14'd10397:data <=32'h0017000D;
14'd10398:data <=32'h0011FFF7;14'd10399:data <=32'h0006FFE6;14'd10400:data <=32'hFFF8FFDB;
14'd10401:data <=32'hFFE8FFD6;14'd10402:data <=32'hFFD9FFD4;14'd10403:data <=32'hFFCBFFD5;
14'd10404:data <=32'hFFBDFFDA;14'd10405:data <=32'hFFB0FFE3;14'd10406:data <=32'hFFA4FFEE;
14'd10407:data <=32'hFF9BFFFC;14'd10408:data <=32'hFF96000C;14'd10409:data <=32'hFF96001D;
14'd10410:data <=32'hFF9A002D;14'd10411:data <=32'hFF9F0039;14'd10412:data <=32'hFFA50044;
14'd10413:data <=32'hFFAA004C;14'd10414:data <=32'hFFAE0055;14'd10415:data <=32'hFFB10060;
14'd10416:data <=32'hFFB6006E;14'd10417:data <=32'hFFBF007F;14'd10418:data <=32'hFFCD008F;
14'd10419:data <=32'hFFE3009E;14'd10420:data <=32'hFFFD00A7;14'd10421:data <=32'h001B00A8;
14'd10422:data <=32'h003600A0;14'd10423:data <=32'h004F0092;14'd10424:data <=32'h0060007F;
14'd10425:data <=32'h006A006A;14'd10426:data <=32'h006F0058;14'd10427:data <=32'h00710049;
14'd10428:data <=32'h0071003C;14'd10429:data <=32'h00700032;14'd10430:data <=32'h006E0028;
14'd10431:data <=32'h006D0022;14'd10432:data <=32'h00DD0091;14'd10433:data <=32'h01070068;
14'd10434:data <=32'h010A0032;14'd10435:data <=32'h0077001C;14'd10436:data <=32'h00510049;
14'd10437:data <=32'h00680050;14'd10438:data <=32'h0086004E;14'd10439:data <=32'h00A70041;
14'd10440:data <=32'h00C50026;14'd10441:data <=32'h00DAFFFF;14'd10442:data <=32'h00E3FFD0;
14'd10443:data <=32'h00DDFF9F;14'd10444:data <=32'h00CAFF72;14'd10445:data <=32'h00AAFF4D;
14'd10446:data <=32'h0085FF30;14'd10447:data <=32'h005BFF1D;14'd10448:data <=32'h002FFF13;
14'd10449:data <=32'h0003FF14;14'd10450:data <=32'hFFD6FF1D;14'd10451:data <=32'hFFAEFF31;
14'd10452:data <=32'hFF8BFF4E;14'd10453:data <=32'hFF72FF73;14'd10454:data <=32'hFF64FF9C;
14'd10455:data <=32'hFF64FFC6;14'd10456:data <=32'hFF6FFFEA;14'd10457:data <=32'hFF830006;
14'd10458:data <=32'hFF9B0019;14'd10459:data <=32'hFFB40023;14'd10460:data <=32'hFFC90023;
14'd10461:data <=32'hFFDA0020;14'd10462:data <=32'hFFE7001B;14'd10463:data <=32'hFFF30015;
14'd10464:data <=32'hFFFB000E;14'd10465:data <=32'h00040005;14'd10466:data <=32'h000CFFFA;
14'd10467:data <=32'h0010FFEC;14'd10468:data <=32'h0011FFDB;14'd10469:data <=32'h000CFFC9;
14'd10470:data <=32'h0001FFB8;14'd10471:data <=32'hFFEFFFA9;14'd10472:data <=32'hFFDAFFA0;
14'd10473:data <=32'hFFC2FF9E;14'd10474:data <=32'hFFA9FFA0;14'd10475:data <=32'hFF8FFFA9;
14'd10476:data <=32'hFF78FFB6;14'd10477:data <=32'hFF62FFC9;14'd10478:data <=32'hFF4EFFE2;
14'd10479:data <=32'hFF3D0001;14'd10480:data <=32'hFF340025;14'd10481:data <=32'hFF320050;
14'd10482:data <=32'hFF3E007C;14'd10483:data <=32'hFF5500A5;14'd10484:data <=32'hFF7A00C8;
14'd10485:data <=32'hFFA700DE;14'd10486:data <=32'hFFD600E6;14'd10487:data <=32'h000500E1;
14'd10488:data <=32'h002C00CF;14'd10489:data <=32'h004B00B5;14'd10490:data <=32'h005E0097;
14'd10491:data <=32'h0068007C;14'd10492:data <=32'h006B0062;14'd10493:data <=32'h0068004C;
14'd10494:data <=32'h0060003A;14'd10495:data <=32'h0057002D;14'd10496:data <=32'h00320097;
14'd10497:data <=32'h004F009C;14'd10498:data <=32'h00710087;14'd10499:data <=32'h006F002D;
14'd10500:data <=32'h003A0052;14'd10501:data <=32'h0043005C;14'd10502:data <=32'h00530062;
14'd10503:data <=32'h00690064;14'd10504:data <=32'h0083005C;14'd10505:data <=32'h009A0049;
14'd10506:data <=32'h00AC002F;14'd10507:data <=32'h00B4000F;14'd10508:data <=32'h00B3FFF0;
14'd10509:data <=32'h00ABFFD3;14'd10510:data <=32'h009EFFBC;14'd10511:data <=32'h008FFFA8;
14'd10512:data <=32'h007EFF99;14'd10513:data <=32'h006CFF8B;14'd10514:data <=32'h0058FF81;
14'd10515:data <=32'h0043FF7A;14'd10516:data <=32'h002CFF77;14'd10517:data <=32'h0017FF79;
14'd10518:data <=32'h0003FF81;14'd10519:data <=32'hFFF4FF8C;14'd10520:data <=32'hFFEAFF9A;
14'd10521:data <=32'hFFE5FFA4;14'd10522:data <=32'hFFE1FFAC;14'd10523:data <=32'hFFDEFFB1;
14'd10524:data <=32'hFFD8FFB6;14'd10525:data <=32'hFFD0FFBC;14'd10526:data <=32'hFFC9FFC6;
14'd10527:data <=32'hFFC2FFD3;14'd10528:data <=32'hFFC1FFE4;14'd10529:data <=32'hFFC7FFF7;
14'd10530:data <=32'hFFD40006;14'd10531:data <=32'hFFE6000E;14'd10532:data <=32'hFFFC0010;
14'd10533:data <=32'h0010000A;14'd10534:data <=32'h0022FFF9;14'd10535:data <=32'h002DFFE5;
14'd10536:data <=32'h0031FFCD;14'd10537:data <=32'h002CFFB2;14'd10538:data <=32'h0021FF9B;
14'd10539:data <=32'h000EFF84;14'd10540:data <=32'hFFF6FF72;14'd10541:data <=32'hFFD5FF65;
14'd10542:data <=32'hFFB0FF5F;14'd10543:data <=32'hFF89FF64;14'd10544:data <=32'hFF61FF76;
14'd10545:data <=32'hFF3BFF92;14'd10546:data <=32'hFF1FFFBB;14'd10547:data <=32'hFF0EFFEB;
14'd10548:data <=32'hFF0C001E;14'd10549:data <=32'hFF18004E;14'd10550:data <=32'hFF300077;
14'd10551:data <=32'hFF4F0095;14'd10552:data <=32'hFF7100A8;14'd10553:data <=32'hFF9300B2;
14'd10554:data <=32'hFFB000B5;14'd10555:data <=32'hFFC900B5;14'd10556:data <=32'hFFE000B2;
14'd10557:data <=32'hFFF400AE;14'd10558:data <=32'h000700A8;14'd10559:data <=32'h001800A0;
14'd10560:data <=32'h0020005E;14'd10561:data <=32'h001F005D;14'd10562:data <=32'h0025006A;
14'd10563:data <=32'h004400B1;14'd10564:data <=32'h002900CA;14'd10565:data <=32'h004500C5;
14'd10566:data <=32'h006300BD;14'd10567:data <=32'h008100AC;14'd10568:data <=32'h009D0095;
14'd10569:data <=32'h00B40074;14'd10570:data <=32'h00C2004C;14'd10571:data <=32'h00C20023;
14'd10572:data <=32'h00B8FFFE;14'd10573:data <=32'h00A3FFE0;14'd10574:data <=32'h0089FFCC;
14'd10575:data <=32'h006FFFC2;14'd10576:data <=32'h0058FFC0;14'd10577:data <=32'h0046FFC4;
14'd10578:data <=32'h0039FFCB;14'd10579:data <=32'h002FFFD2;14'd10580:data <=32'h002AFFDA;
14'd10581:data <=32'h0028FFE1;14'd10582:data <=32'h0029FFE8;14'd10583:data <=32'h002EFFED;
14'd10584:data <=32'h0036FFEF;14'd10585:data <=32'h0040FFEC;14'd10586:data <=32'h0049FFE3;
14'd10587:data <=32'h004EFFD4;14'd10588:data <=32'h004CFFC1;14'd10589:data <=32'h0043FFAF;
14'd10590:data <=32'h0032FFA2;14'd10591:data <=32'h001CFF9C;14'd10592:data <=32'h0007FF9E;
14'd10593:data <=32'hFFF4FFA9;14'd10594:data <=32'hFFE7FFB9;14'd10595:data <=32'hFFE4FFCA;
14'd10596:data <=32'hFFE8FFDB;14'd10597:data <=32'hFFF0FFE7;14'd10598:data <=32'hFFFCFFED;
14'd10599:data <=32'h0008FFED;14'd10600:data <=32'h0014FFE9;14'd10601:data <=32'h001DFFE1;
14'd10602:data <=32'h0024FFD6;14'd10603:data <=32'h0029FFC8;14'd10604:data <=32'h002AFFB7;
14'd10605:data <=32'h0026FFA4;14'd10606:data <=32'h001CFF91;14'd10607:data <=32'h000BFF80;
14'd10608:data <=32'hFFF4FF73;14'd10609:data <=32'hFFD7FF6C;14'd10610:data <=32'hFFBBFF6D;
14'd10611:data <=32'hFF9FFF76;14'd10612:data <=32'hFF88FF86;14'd10613:data <=32'hFF77FF99;
14'd10614:data <=32'hFF6AFFAC;14'd10615:data <=32'hFF63FFBE;14'd10616:data <=32'hFF5CFFCD;
14'd10617:data <=32'hFF54FFDB;14'd10618:data <=32'hFF49FFEB;14'd10619:data <=32'hFF3D0000;
14'd10620:data <=32'hFF330019;14'd10621:data <=32'hFF2C0039;14'd10622:data <=32'hFF2F005C;
14'd10623:data <=32'hFF390082;14'd10624:data <=32'hFFE60086;14'd10625:data <=32'hFFEC007F;
14'd10626:data <=32'hFFDD007A;14'd10627:data <=32'hFF6300B6;14'd10628:data <=32'hFF5200F6;
14'd10629:data <=32'hFF810117;14'd10630:data <=32'hFFB9012B;14'd10631:data <=32'hFFF50134;
14'd10632:data <=32'h0034012B;14'd10633:data <=32'h006F0113;14'd10634:data <=32'h00A000EA;
14'd10635:data <=32'h00C300B7;14'd10636:data <=32'h00D3007F;14'd10637:data <=32'h00D40049;
14'd10638:data <=32'h00C5001A;14'd10639:data <=32'h00AEFFF6;14'd10640:data <=32'h0091FFDD;
14'd10641:data <=32'h0073FFCF;14'd10642:data <=32'h0059FFCB;14'd10643:data <=32'h0041FFCB;
14'd10644:data <=32'h002CFFD0;14'd10645:data <=32'h001CFFDB;14'd10646:data <=32'h0011FFE9;
14'd10647:data <=32'h000BFFF9;14'd10648:data <=32'h000D000A;14'd10649:data <=32'h00160018;
14'd10650:data <=32'h0024001F;14'd10651:data <=32'h00350020;14'd10652:data <=32'h00430019;
14'd10653:data <=32'h004E000D;14'd10654:data <=32'h0052FFFE;14'd10655:data <=32'h0051FFF1;
14'd10656:data <=32'h004CFFE6;14'd10657:data <=32'h0045FFE1;14'd10658:data <=32'h003EFFDE;
14'd10659:data <=32'h003CFFDE;14'd10660:data <=32'h003CFFDD;14'd10661:data <=32'h003EFFD9;
14'd10662:data <=32'h003FFFD3;14'd10663:data <=32'h003FFFCA;14'd10664:data <=32'h003BFFC1;
14'd10665:data <=32'h0034FFB8;14'd10666:data <=32'h002CFFB3;14'd10667:data <=32'h0023FFB0;
14'd10668:data <=32'h001BFFAD;14'd10669:data <=32'h0015FFAD;14'd10670:data <=32'h000EFFAE;
14'd10671:data <=32'h0009FFAE;14'd10672:data <=32'h0004FFAE;14'd10673:data <=32'hFFFFFFAD;
14'd10674:data <=32'hFFFAFFAF;14'd10675:data <=32'hFFF8FFB1;14'd10676:data <=32'hFFF8FFB2;
14'd10677:data <=32'hFFFAFFB1;14'd10678:data <=32'hFFFDFFAA;14'd10679:data <=32'h0000FF9F;
14'd10680:data <=32'hFFFDFF8C;14'd10681:data <=32'hFFF0FF75;14'd10682:data <=32'hFFD8FF60;
14'd10683:data <=32'hFFB6FF51;14'd10684:data <=32'hFF8BFF4D;14'd10685:data <=32'hFF5DFF58;
14'd10686:data <=32'hFF30FF6F;14'd10687:data <=32'hFF0CFF94;14'd10688:data <=32'hFF650015;
14'd10689:data <=32'hFF5B0021;14'd10690:data <=32'hFF560019;14'd10691:data <=32'hFF15FFD7;
14'd10692:data <=32'hFED90025;14'd10693:data <=32'hFEE2005E;14'd10694:data <=32'hFEF80095;
14'd10695:data <=32'hFF1B00C5;14'd10696:data <=32'hFF4B00EC;14'd10697:data <=32'hFF820104;
14'd10698:data <=32'hFFBD010B;14'd10699:data <=32'hFFF20102;14'd10700:data <=32'h002000ED;
14'd10701:data <=32'h004300D0;14'd10702:data <=32'h005A00B1;14'd10703:data <=32'h00670093;
14'd10704:data <=32'h006D0077;14'd10705:data <=32'h006F0061;14'd10706:data <=32'h0071004B;
14'd10707:data <=32'h006F0038;14'd10708:data <=32'h006A0025;14'd10709:data <=32'h00620015;
14'd10710:data <=32'h00580007;14'd10711:data <=32'h004AFFFD;14'd10712:data <=32'h003DFFF9;
14'd10713:data <=32'h0032FFFA;14'd10714:data <=32'h002AFFFC;14'd10715:data <=32'h0024FFFF;
14'd10716:data <=32'h00200002;14'd10717:data <=32'h001D0004;14'd10718:data <=32'h00170007;
14'd10719:data <=32'h0012000B;14'd10720:data <=32'h000F0013;14'd10721:data <=32'h000D001F;
14'd10722:data <=32'h0012002C;14'd10723:data <=32'h001F0039;14'd10724:data <=32'h00310042;
14'd10725:data <=32'h00480042;14'd10726:data <=32'h0060003B;14'd10727:data <=32'h0074002B;
14'd10728:data <=32'h00830014;14'd10729:data <=32'h008AFFF9;14'd10730:data <=32'h0089FFDE;
14'd10731:data <=32'h0080FFC6;14'd10732:data <=32'h0073FFB2;14'd10733:data <=32'h0062FFA3;
14'd10734:data <=32'h004FFF99;14'd10735:data <=32'h003EFF94;14'd10736:data <=32'h002BFF92;
14'd10737:data <=32'h001AFF96;14'd10738:data <=32'h000BFF9E;14'd10739:data <=32'h0001FFA9;
14'd10740:data <=32'hFFFEFFB7;14'd10741:data <=32'h0002FFC3;14'd10742:data <=32'h000DFFCA;
14'd10743:data <=32'h001CFFCA;14'd10744:data <=32'h002CFFBF;14'd10745:data <=32'h0036FFA9;
14'd10746:data <=32'h0037FF8E;14'd10747:data <=32'h002BFF6F;14'd10748:data <=32'h0014FF53;
14'd10749:data <=32'hFFF3FF40;14'd10750:data <=32'hFFCAFF37;14'd10751:data <=32'hFFA0FF39;
14'd10752:data <=32'hFFC6FF55;14'd10753:data <=32'hFF9AFF47;14'd10754:data <=32'hFF81FF4A;
14'd10755:data <=32'hFF96FF71;14'd10756:data <=32'hFF4BFF9F;14'd10757:data <=32'hFF3FFFBC;
14'd10758:data <=32'hFF37FFDA;14'd10759:data <=32'hFF36FFFA;14'd10760:data <=32'hFF3D001A;
14'd10761:data <=32'hFF4A0035;14'd10762:data <=32'hFF5D004A;14'd10763:data <=32'hFF700058;
14'd10764:data <=32'hFF81005F;14'd10765:data <=32'hFF8F0064;14'd10766:data <=32'hFF98006A;
14'd10767:data <=32'hFF9F0072;14'd10768:data <=32'hFFA7007D;14'd10769:data <=32'hFFB5008C;
14'd10770:data <=32'hFFC80098;14'd10771:data <=32'hFFE000A1;14'd10772:data <=32'hFFFB00A4;
14'd10773:data <=32'h0018009F;14'd10774:data <=32'h00320092;14'd10775:data <=32'h00460081;
14'd10776:data <=32'h0055006A;14'd10777:data <=32'h005F0054;14'd10778:data <=32'h0063003D;
14'd10779:data <=32'h00630025;14'd10780:data <=32'h005D000F;14'd10781:data <=32'h0051FFFA;
14'd10782:data <=32'h003EFFE9;14'd10783:data <=32'h0027FFDF;14'd10784:data <=32'h000DFFDF;
14'd10785:data <=32'hFFF3FFE9;14'd10786:data <=32'hFFE0FFFC;14'd10787:data <=32'hFFD40017;
14'd10788:data <=32'hFFD50034;14'd10789:data <=32'hFFE1004F;14'd10790:data <=32'hFFF60064;
14'd10791:data <=32'h00110071;14'd10792:data <=32'h002E0073;14'd10793:data <=32'h0049006E;
14'd10794:data <=32'h00600062;14'd10795:data <=32'h00730051;14'd10796:data <=32'h0081003F;
14'd10797:data <=32'h008A002B;14'd10798:data <=32'h00910017;14'd10799:data <=32'h00930003;
14'd10800:data <=32'h0092FFED;14'd10801:data <=32'h008DFFD9;14'd10802:data <=32'h0085FFC8;
14'd10803:data <=32'h007AFFBA;14'd10804:data <=32'h006FFFB1;14'd10805:data <=32'h0066FFAB;
14'd10806:data <=32'h005FFFA6;14'd10807:data <=32'h005CFFA0;14'd10808:data <=32'h005AFF96;
14'd10809:data <=32'h0057FF87;14'd10810:data <=32'h0050FF74;14'd10811:data <=32'h0040FF61;
14'd10812:data <=32'h002AFF4F;14'd10813:data <=32'h000DFF44;14'd10814:data <=32'hFFEDFF42;
14'd10815:data <=32'hFFCDFF48;14'd10816:data <=32'h0078FF7D;14'd10817:data <=32'h0067FF45;
14'd10818:data <=32'h003AFF25;14'd10819:data <=32'hFFBBFF79;14'd10820:data <=32'hFF7FFFA5;
14'd10821:data <=32'hFF81FFBD;14'd10822:data <=32'hFF87FFD0;14'd10823:data <=32'hFF90FFDF;
14'd10824:data <=32'hFF9BFFEB;14'd10825:data <=32'hFFA8FFF1;14'd10826:data <=32'hFFB5FFF0;
14'd10827:data <=32'hFFBDFFEA;14'd10828:data <=32'hFFBEFFDF;14'd10829:data <=32'hFFB7FFD4;
14'd10830:data <=32'hFFA6FFCD;14'd10831:data <=32'hFF90FFCD;14'd10832:data <=32'hFF77FFDA;
14'd10833:data <=32'hFF64FFF2;14'd10834:data <=32'hFF580011;14'd10835:data <=32'hFF570033;
14'd10836:data <=32'hFF620055;14'd10837:data <=32'hFF760072;14'd10838:data <=32'hFF900088;
14'd10839:data <=32'hFFAD0097;14'd10840:data <=32'hFFCB009D;14'd10841:data <=32'hFFEA009D;
14'd10842:data <=32'h00080096;14'd10843:data <=32'h0022008A;14'd10844:data <=32'h00390076;
14'd10845:data <=32'h0048005D;14'd10846:data <=32'h00500040;14'd10847:data <=32'h004E0023;
14'd10848:data <=32'h0043000A;14'd10849:data <=32'h002FFFF8;14'd10850:data <=32'h0018FFEF;
14'd10851:data <=32'h0001FFF0;14'd10852:data <=32'hFFEDFFF9;14'd10853:data <=32'hFFDF0008;
14'd10854:data <=32'hFFD80019;14'd10855:data <=32'hFFD70029;14'd10856:data <=32'hFFDA0037;
14'd10857:data <=32'hFFDF0044;14'd10858:data <=32'hFFE4004F;14'd10859:data <=32'hFFEC005C;
14'd10860:data <=32'hFFF40067;14'd10861:data <=32'h00000074;14'd10862:data <=32'h00120080;
14'd10863:data <=32'h0027008A;14'd10864:data <=32'h0041008F;14'd10865:data <=32'h005F008D;
14'd10866:data <=32'h007B0085;14'd10867:data <=32'h00960077;14'd10868:data <=32'h00AF0063;
14'd10869:data <=32'h00C6004B;14'd10870:data <=32'h00D9002E;14'd10871:data <=32'h00E9000D;
14'd10872:data <=32'h00F3FFE5;14'd10873:data <=32'h00F6FFB9;14'd10874:data <=32'h00EDFF87;
14'd10875:data <=32'h00D9FF58;14'd10876:data <=32'h00B5FF2D;14'd10877:data <=32'h0087FF0E;
14'd10878:data <=32'h0051FEFC;14'd10879:data <=32'h001AFEFA;14'd10880:data <=32'h007BFFD5;
14'd10881:data <=32'h008BFFAC;14'd10882:data <=32'h0084FF72;14'd10883:data <=32'hFFFBFF1D;
14'd10884:data <=32'hFFA6FF4B;14'd10885:data <=32'hFF97FF6C;14'd10886:data <=32'hFF8FFF8B;
14'd10887:data <=32'hFF90FFA8;14'd10888:data <=32'hFF97FFC2;14'd10889:data <=32'hFFA3FFD6;
14'd10890:data <=32'hFFB6FFE2;14'd10891:data <=32'hFFC8FFE5;14'd10892:data <=32'hFFD7FFDF;
14'd10893:data <=32'hFFDFFFD2;14'd10894:data <=32'hFFDDFFC2;14'd10895:data <=32'hFFD1FFB5;
14'd10896:data <=32'hFFBEFFAD;14'd10897:data <=32'hFFA8FFB1;14'd10898:data <=32'hFF94FFBC;
14'd10899:data <=32'hFF85FFCE;14'd10900:data <=32'hFF7DFFE5;14'd10901:data <=32'hFF7BFFFA;
14'd10902:data <=32'hFF7E000E;14'd10903:data <=32'hFF85001F;14'd10904:data <=32'hFF8E002E;
14'd10905:data <=32'hFF98003B;14'd10906:data <=32'hFFA40046;14'd10907:data <=32'hFFB20050;
14'd10908:data <=32'hFFC20056;14'd10909:data <=32'hFFD40058;14'd10910:data <=32'hFFE40055;
14'd10911:data <=32'hFFF1004E;14'd10912:data <=32'hFFFA0044;14'd10913:data <=32'hFFFE003A;
14'd10914:data <=32'h00000032;14'd10915:data <=32'hFFFF002C;14'd10916:data <=32'hFFFC0029;
14'd10917:data <=32'hFFFD0026;14'd10918:data <=32'hFFFF0023;14'd10919:data <=32'h0000001E;
14'd10920:data <=32'hFFFE0017;14'd10921:data <=32'hFFF8000E;14'd10922:data <=32'hFFED0008;
14'd10923:data <=32'hFFDD0005;14'd10924:data <=32'hFFCA000A;14'd10925:data <=32'hFFB70019;
14'd10926:data <=32'hFFA90030;14'd10927:data <=32'hFFA2004D;14'd10928:data <=32'hFFA4006E;
14'd10929:data <=32'hFFB10090;14'd10930:data <=32'hFFC800AE;14'd10931:data <=32'hFFE800C8;
14'd10932:data <=32'h000E00DA;14'd10933:data <=32'h003A00E3;14'd10934:data <=32'h006900E4;
14'd10935:data <=32'h009C00D9;14'd10936:data <=32'h00CE00C1;14'd10937:data <=32'h00FC009C;
14'd10938:data <=32'h011F006A;14'd10939:data <=32'h0137002C;14'd10940:data <=32'h013BFFEA;
14'd10941:data <=32'h012DFFA9;14'd10942:data <=32'h010EFF70;14'd10943:data <=32'h00E3FF44;
14'd10944:data <=32'h00A0FFC6;14'd10945:data <=32'h00A8FFA9;14'd10946:data <=32'h00B9FF88;
14'd10947:data <=32'h00CDFF4C;14'd10948:data <=32'h0073FF50;14'd10949:data <=32'h0058FF4B;
14'd10950:data <=32'h003EFF4B;14'd10951:data <=32'h0026FF4C;14'd10952:data <=32'h000FFF52;
14'd10953:data <=32'hFFFAFF5B;14'd10954:data <=32'hFFEBFF67;14'd10955:data <=32'hFFE0FF71;
14'd10956:data <=32'hFFD8FF7A;14'd10957:data <=32'hFFCEFF7F;14'd10958:data <=32'hFFC3FF83;
14'd10959:data <=32'hFFB6FF8A;14'd10960:data <=32'hFFA6FF94;14'd10961:data <=32'hFF96FFA3;
14'd10962:data <=32'hFF8DFFB9;14'd10963:data <=32'hFF89FFD0;14'd10964:data <=32'hFF8DFFE9;
14'd10965:data <=32'hFF98FFFC;14'd10966:data <=32'hFFA8000A;14'd10967:data <=32'hFFB8000F;
14'd10968:data <=32'hFFC7000E;14'd10969:data <=32'hFFD10009;14'd10970:data <=32'hFFD60003;
14'd10971:data <=32'hFFD8FFFD;14'd10972:data <=32'hFFD6FFF8;14'd10973:data <=32'hFFD3FFF5;
14'd10974:data <=32'hFFCFFFF2;14'd10975:data <=32'hFFC9FFF2;14'd10976:data <=32'hFFC2FFF4;
14'd10977:data <=32'hFFBCFFF7;14'd10978:data <=32'hFFB4FFFF;14'd10979:data <=32'hFFAF000B;
14'd10980:data <=32'hFFAE0019;14'd10981:data <=32'hFFB30027;14'd10982:data <=32'hFFBD0034;
14'd10983:data <=32'hFFCC003A;14'd10984:data <=32'hFFDC0039;14'd10985:data <=32'hFFEA0031;
14'd10986:data <=32'hFFF10025;14'd10987:data <=32'hFFF10015;14'd10988:data <=32'hFFE70008;
14'd10989:data <=32'hFFD70000;14'd10990:data <=32'hFFC30001;14'd10991:data <=32'hFFAF000A;
14'd10992:data <=32'hFF9F001B;14'd10993:data <=32'hFF940033;14'd10994:data <=32'hFF91004D;
14'd10995:data <=32'hFF940069;14'd10996:data <=32'hFF9E0086;14'd10997:data <=32'hFFAE00A2;
14'd10998:data <=32'hFFC700BC;14'd10999:data <=32'hFFE600D1;14'd11000:data <=32'h000D00DF;
14'd11001:data <=32'h003800E3;14'd11002:data <=32'h006600DC;14'd11003:data <=32'h009100C8;
14'd11004:data <=32'h00B400AA;14'd11005:data <=32'h00CD0084;14'd11006:data <=32'h00DB005D;
14'd11007:data <=32'h00DF0037;14'd11008:data <=32'h00F90045;14'd11009:data <=32'h0110001B;
14'd11010:data <=32'h01140001;14'd11011:data <=32'h00E4003E;14'd11012:data <=32'h00B90038;
14'd11013:data <=32'h00C80023;14'd11014:data <=32'h00D50006;14'd11015:data <=32'h00DCFFE5;
14'd11016:data <=32'h00DBFFC0;14'd11017:data <=32'h00D3FF9D;14'd11018:data <=32'h00C2FF7C;
14'd11019:data <=32'h00ABFF5E;14'd11020:data <=32'h0090FF43;14'd11021:data <=32'h006FFF2C;
14'd11022:data <=32'h0048FF1B;14'd11023:data <=32'h001BFF12;14'd11024:data <=32'hFFECFF14;
14'd11025:data <=32'hFFBDFF24;14'd11026:data <=32'hFF94FF42;14'd11027:data <=32'hFF77FF69;
14'd11028:data <=32'hFF67FF96;14'd11029:data <=32'hFF67FFC2;14'd11030:data <=32'hFF74FFEA;
14'd11031:data <=32'hFF8A0008;14'd11032:data <=32'hFFA5001A;14'd11033:data <=32'hFFC10023;
14'd11034:data <=32'hFFD80022;14'd11035:data <=32'hFFEE001C;14'd11036:data <=32'hFFFE0011;
14'd11037:data <=32'h00090003;14'd11038:data <=32'h0010FFF2;14'd11039:data <=32'h0010FFE1;
14'd11040:data <=32'h000CFFD0;14'd11041:data <=32'h0000FFC1;14'd11042:data <=32'hFFF0FFB5;
14'd11043:data <=32'hFFDEFFB1;14'd11044:data <=32'hFFC9FFB5;14'd11045:data <=32'hFFB9FFBE;
14'd11046:data <=32'hFFADFFCA;14'd11047:data <=32'hFFA6FFD9;14'd11048:data <=32'hFFA6FFE6;
14'd11049:data <=32'hFFA8FFED;14'd11050:data <=32'hFFA9FFF4;14'd11051:data <=32'hFFA8FFF5;
14'd11052:data <=32'hFFA4FFF9;14'd11053:data <=32'hFF9CFFFC;14'd11054:data <=32'hFF930005;
14'd11055:data <=32'hFF8B0013;14'd11056:data <=32'hFF870023;14'd11057:data <=32'hFF870037;
14'd11058:data <=32'hFF8C0049;14'd11059:data <=32'hFF96005A;14'd11060:data <=32'hFFA20069;
14'd11061:data <=32'hFFAF0074;14'd11062:data <=32'hFFBD007D;14'd11063:data <=32'hFFCC0085;
14'd11064:data <=32'hFFDC008B;14'd11065:data <=32'hFFED008F;14'd11066:data <=32'hFFFF008F;
14'd11067:data <=32'h0011008A;14'd11068:data <=32'h001E0083;14'd11069:data <=32'h00280079;
14'd11070:data <=32'h002C0072;14'd11071:data <=32'h002C006E;14'd11072:data <=32'h007100EA;
14'd11073:data <=32'h00A100DF;14'd11074:data <=32'h00B700BF;14'd11075:data <=32'h003B008B;
14'd11076:data <=32'h001700A7;14'd11077:data <=32'h003900B5;14'd11078:data <=32'h006100B9;
14'd11079:data <=32'h008C00AF;14'd11080:data <=32'h00B3009A;14'd11081:data <=32'h00D5007B;
14'd11082:data <=32'h00EE0055;14'd11083:data <=32'h01000029;14'd11084:data <=32'h0108FFFA;
14'd11085:data <=32'h0105FFC7;14'd11086:data <=32'h00F7FF94;14'd11087:data <=32'h00DAFF65;
14'd11088:data <=32'h00B2FF3E;14'd11089:data <=32'h0081FF23;14'd11090:data <=32'h004BFF19;
14'd11091:data <=32'h0016FF1F;14'd11092:data <=32'hFFE7FF33;14'd11093:data <=32'hFFC5FF50;
14'd11094:data <=32'hFFAFFF73;14'd11095:data <=32'hFFA4FF95;14'd11096:data <=32'hFFA3FFB3;
14'd11097:data <=32'hFFA7FFCD;14'd11098:data <=32'hFFB0FFE3;14'd11099:data <=32'hFFBBFFF3;
14'd11100:data <=32'hFFC90000;14'd11101:data <=32'hFFD8000B;14'd11102:data <=32'hFFEA000F;
14'd11103:data <=32'hFFFC0010;14'd11104:data <=32'h000C000A;14'd11105:data <=32'h001BFFFF;
14'd11106:data <=32'h0025FFF1;14'd11107:data <=32'h0029FFE0;14'd11108:data <=32'h0028FFCF;
14'd11109:data <=32'h0024FFBF;14'd11110:data <=32'h001CFFB1;14'd11111:data <=32'h0013FFA6;
14'd11112:data <=32'h0009FF9A;14'd11113:data <=32'hFFFBFF8F;14'd11114:data <=32'hFFEAFF82;
14'd11115:data <=32'hFFD4FF79;14'd11116:data <=32'hFFB8FF74;14'd11117:data <=32'hFF98FF77;
14'd11118:data <=32'hFF75FF85;14'd11119:data <=32'hFF57FF9C;14'd11120:data <=32'hFF3EFFBC;
14'd11121:data <=32'hFF30FFE3;14'd11122:data <=32'hFF2E000D;14'd11123:data <=32'hFF370034;
14'd11124:data <=32'hFF480057;14'd11125:data <=32'hFF600072;14'd11126:data <=32'hFF7C0085;
14'd11127:data <=32'hFF980091;14'd11128:data <=32'hFFB50096;14'd11129:data <=32'hFFD10094;
14'd11130:data <=32'hFFEA008D;14'd11131:data <=32'hFFFD0080;14'd11132:data <=32'h000B006D;
14'd11133:data <=32'h00110059;14'd11134:data <=32'h000C0048;14'd11135:data <=32'hFFFF003C;
14'd11136:data <=32'hFFC00099;14'd11137:data <=32'hFFCE00B1;14'd11138:data <=32'hFFF000B5;
14'd11139:data <=32'h00080063;14'd11140:data <=32'hFFCF007D;14'd11141:data <=32'hFFDF0093;
14'd11142:data <=32'hFFF500A5;14'd11143:data <=32'h001300AF;14'd11144:data <=32'h003200B3;
14'd11145:data <=32'h005100AC;14'd11146:data <=32'h006C00A0;14'd11147:data <=32'h00870090;
14'd11148:data <=32'h009E007A;14'd11149:data <=32'h00B20060;14'd11150:data <=32'h00C00040;
14'd11151:data <=32'h00C6001D;14'd11152:data <=32'h00C4FFF8;14'd11153:data <=32'h00B8FFD7;
14'd11154:data <=32'h00A4FFBC;14'd11155:data <=32'h008AFFA8;14'd11156:data <=32'h0071FF9E;
14'd11157:data <=32'h005AFF9C;14'd11158:data <=32'h0048FF9C;14'd11159:data <=32'h003BFF9E;
14'd11160:data <=32'h0030FF9F;14'd11161:data <=32'h0025FF9F;14'd11162:data <=32'h0019FF9E;
14'd11163:data <=32'h000AFFA0;14'd11164:data <=32'hFFFBFFA5;14'd11165:data <=32'hFFEDFFB0;
14'd11166:data <=32'hFFE2FFBE;14'd11167:data <=32'hFFDCFFD0;14'd11168:data <=32'hFFDEFFE2;
14'd11169:data <=32'hFFE3FFF2;14'd11170:data <=32'hFFEEFFFF;14'd11171:data <=32'hFFFC0007;
14'd11172:data <=32'h000C000B;14'd11173:data <=32'h001D000C;14'd11174:data <=32'h00300007;
14'd11175:data <=32'h0041FFFD;14'd11176:data <=32'h0052FFEB;14'd11177:data <=32'h005FFFD4;
14'd11178:data <=32'h0065FFB4;14'd11179:data <=32'h0060FF91;14'd11180:data <=32'h0051FF6E;
14'd11181:data <=32'h0035FF4D;14'd11182:data <=32'h000EFF36;14'd11183:data <=32'hFFE0FF2B;
14'd11184:data <=32'hFFB0FF2F;14'd11185:data <=32'hFF83FF40;14'd11186:data <=32'hFF5DFF5C;
14'd11187:data <=32'hFF42FF7F;14'd11188:data <=32'hFF31FFA6;14'd11189:data <=32'hFF2AFFCC;
14'd11190:data <=32'hFF2AFFF1;14'd11191:data <=32'hFF320012;14'd11192:data <=32'hFF3E002F;
14'd11193:data <=32'hFF4F004A;14'd11194:data <=32'hFF65005E;14'd11195:data <=32'hFF7C006A;
14'd11196:data <=32'hFF940071;14'd11197:data <=32'hFFA90070;14'd11198:data <=32'hFFB7006B;
14'd11199:data <=32'hFFBF0065;14'd11200:data <=32'hFFD6002E;14'd11201:data <=32'hFFC3002F;
14'd11202:data <=32'hFFB90045;14'd11203:data <=32'hFFC60097;14'd11204:data <=32'hFF9E00AE;
14'd11205:data <=32'hFFBA00BF;14'd11206:data <=32'hFFDC00C8;14'd11207:data <=32'h000100C9;
14'd11208:data <=32'h002200C0;14'd11209:data <=32'h003E00AE;14'd11210:data <=32'h00530099;
14'd11211:data <=32'h00610081;14'd11212:data <=32'h0069006A;14'd11213:data <=32'h006D0056;
14'd11214:data <=32'h006E0042;14'd11215:data <=32'h006C0031;14'd11216:data <=32'h00650021;
14'd11217:data <=32'h005C0014;14'd11218:data <=32'h004F000C;14'd11219:data <=32'h0044000B;
14'd11220:data <=32'h003A000F;14'd11221:data <=32'h00380017;14'd11222:data <=32'h003C001F;
14'd11223:data <=32'h00460024;14'd11224:data <=32'h00550021;14'd11225:data <=32'h00640017;
14'd11226:data <=32'h006E0005;14'd11227:data <=32'h0070FFEF;14'd11228:data <=32'h006AFFDA;
14'd11229:data <=32'h005FFFC8;14'd11230:data <=32'h004CFFBC;14'd11231:data <=32'h003AFFB6;
14'd11232:data <=32'h0027FFB7;14'd11233:data <=32'h0018FFBD;14'd11234:data <=32'h000BFFC5;
14'd11235:data <=32'h0002FFD1;14'd11236:data <=32'hFFFEFFDF;14'd11237:data <=32'hFFFEFFED;
14'd11238:data <=32'h0002FFFC;14'd11239:data <=32'h000E0008;14'd11240:data <=32'h001F000F;
14'd11241:data <=32'h00350011;14'd11242:data <=32'h004B000A;14'd11243:data <=32'h0060FFFA;
14'd11244:data <=32'h006EFFE0;14'd11245:data <=32'h0074FFC3;14'd11246:data <=32'h006FFFA3;
14'd11247:data <=32'h0061FF87;14'd11248:data <=32'h004CFF70;14'd11249:data <=32'h0032FF60;
14'd11250:data <=32'h0019FF58;14'd11251:data <=32'h0001FF55;14'd11252:data <=32'hFFEAFF56;
14'd11253:data <=32'hFFD5FF57;14'd11254:data <=32'hFFBFFF59;14'd11255:data <=32'hFFA9FF5E;
14'd11256:data <=32'hFF92FF65;14'd11257:data <=32'hFF7AFF70;14'd11258:data <=32'hFF64FF80;
14'd11259:data <=32'hFF51FF95;14'd11260:data <=32'hFF41FFAC;14'd11261:data <=32'hFF34FFC4;
14'd11262:data <=32'hFF2BFFDE;14'd11263:data <=32'hFF22FFF9;14'd11264:data <=32'hFFC80037;
14'd11265:data <=32'hFFC20027;14'd11266:data <=32'hFFA4001B;14'd11267:data <=32'hFF14003B;
14'd11268:data <=32'hFEE70075;14'd11269:data <=32'hFF0400AC;14'd11270:data <=32'hFF3100D9;
14'd11271:data <=32'hFF6800F9;14'd11272:data <=32'hFFA30105;14'd11273:data <=32'hFFDD0102;
14'd11274:data <=32'h000E00F0;14'd11275:data <=32'h003500D6;14'd11276:data <=32'h005300B7;
14'd11277:data <=32'h00670093;14'd11278:data <=32'h00710071;14'd11279:data <=32'h00730050;
14'd11280:data <=32'h006D0032;14'd11281:data <=32'h005E0018;14'd11282:data <=32'h00490006;
14'd11283:data <=32'h0031FFFD;14'd11284:data <=32'h001AFFFF;14'd11285:data <=32'h0008000A;
14'd11286:data <=32'hFFFE001B;14'd11287:data <=32'hFFFE002F;14'd11288:data <=32'h0008003E;
14'd11289:data <=32'h00160049;14'd11290:data <=32'h0029004B;14'd11291:data <=32'h00380047;
14'd11292:data <=32'h0046003B;14'd11293:data <=32'h004C002E;14'd11294:data <=32'h00500023;
14'd11295:data <=32'h00500019;14'd11296:data <=32'h004E0010;14'd11297:data <=32'h004E0009;
14'd11298:data <=32'h004C0003;14'd11299:data <=32'h004AFFFD;14'd11300:data <=32'h0046FFF7;
14'd11301:data <=32'h0042FFF2;14'd11302:data <=32'h003EFFF0;14'd11303:data <=32'h0039FFF0;
14'd11304:data <=32'h0037FFF1;14'd11305:data <=32'h0038FFF3;14'd11306:data <=32'h003CFFF4;
14'd11307:data <=32'h0040FFF2;14'd11308:data <=32'h0045FFEC;14'd11309:data <=32'h0048FFE4;
14'd11310:data <=32'h0048FFDB;14'd11311:data <=32'h0044FFD5;14'd11312:data <=32'h003FFFD0;
14'd11313:data <=32'h003BFFD0;14'd11314:data <=32'h003CFFD1;14'd11315:data <=32'h0042FFD0;
14'd11316:data <=32'h004BFFCD;14'd11317:data <=32'h0057FFC2;14'd11318:data <=32'h0060FFAF;
14'd11319:data <=32'h0065FF95;14'd11320:data <=32'h0060FF77;14'd11321:data <=32'h0051FF58;
14'd11322:data <=32'h003AFF3A;14'd11323:data <=32'h001AFF22;14'd11324:data <=32'hFFF3FF11;
14'd11325:data <=32'hFFC7FF09;14'd11326:data <=32'hFF98FF08;14'd11327:data <=32'hFF66FF13;
14'd11328:data <=32'hFF94FFC0;14'd11329:data <=32'hFF86FFB7;14'd11330:data <=32'hFF78FFA1;
14'd11331:data <=32'hFF38FF47;14'd11332:data <=32'hFED9FF7D;14'd11333:data <=32'hFEC6FFBE;
14'd11334:data <=32'hFEC6FFFF;14'd11335:data <=32'hFED8003E;14'd11336:data <=32'hFEF80071;
14'd11337:data <=32'hFF200097;14'd11338:data <=32'hFF4B00B0;14'd11339:data <=32'hFF7600BD;
14'd11340:data <=32'hFF9E00C2;14'd11341:data <=32'hFFC300BF;14'd11342:data <=32'hFFE400B6;
14'd11343:data <=32'h000100A8;14'd11344:data <=32'h00180095;14'd11345:data <=32'h002A007F;
14'd11346:data <=32'h00330067;14'd11347:data <=32'h00340051;14'd11348:data <=32'h0030003F;
14'd11349:data <=32'h00270034;14'd11350:data <=32'h001F002E;14'd11351:data <=32'h001A002D;
14'd11352:data <=32'h0018002D;14'd11353:data <=32'h0019002D;14'd11354:data <=32'h001B002A;
14'd11355:data <=32'h001B0024;14'd11356:data <=32'h0017001E;14'd11357:data <=32'h0011001A;
14'd11358:data <=32'h0009001C;14'd11359:data <=32'h00000020;14'd11360:data <=32'hFFFB002B;
14'd11361:data <=32'hFFFC0038;14'd11362:data <=32'h00020045;14'd11363:data <=32'h000E004F;
14'd11364:data <=32'h001D0055;14'd11365:data <=32'h002D0057;14'd11366:data <=32'h003D0052;
14'd11367:data <=32'h004D004C;14'd11368:data <=32'h005A0043;14'd11369:data <=32'h00650037;
14'd11370:data <=32'h006E0027;14'd11371:data <=32'h00740017;14'd11372:data <=32'h00760003;
14'd11373:data <=32'h0073FFF0;14'd11374:data <=32'h0068FFDE;14'd11375:data <=32'h0059FFD2;
14'd11376:data <=32'h0048FFCD;14'd11377:data <=32'h0036FFD0;14'd11378:data <=32'h002AFFDB;
14'd11379:data <=32'h0026FFEB;14'd11380:data <=32'h002CFFFA;14'd11381:data <=32'h003B0005;
14'd11382:data <=32'h00510007;14'd11383:data <=32'h006A0000;14'd11384:data <=32'h007FFFED;
14'd11385:data <=32'h008FFFD2;14'd11386:data <=32'h0097FFB1;14'd11387:data <=32'h0095FF8D;
14'd11388:data <=32'h008BFF69;14'd11389:data <=32'h0077FF46;14'd11390:data <=32'h005BFF27;
14'd11391:data <=32'h0036FF0B;14'd11392:data <=32'h0037FF48;14'd11393:data <=32'h001AFF1E;
14'd11394:data <=32'h0001FF0B;14'd11395:data <=32'h0004FF20;14'd11396:data <=32'hFFA0FF29;
14'd11397:data <=32'hFF7EFF42;14'd11398:data <=32'hFF66FF60;14'd11399:data <=32'hFF55FF82;
14'd11400:data <=32'hFF4FFFA1;14'd11401:data <=32'hFF4FFFBB;14'd11402:data <=32'hFF50FFD0;
14'd11403:data <=32'hFF52FFE1;14'd11404:data <=32'hFF53FFF3;14'd11405:data <=32'hFF530006;
14'd11406:data <=32'hFF56001B;14'd11407:data <=32'hFF5B0032;14'd11408:data <=32'hFF660047;
14'd11409:data <=32'hFF74005A;14'd11410:data <=32'hFF870069;14'd11411:data <=32'hFF990075;
14'd11412:data <=32'hFFAC007D;14'd11413:data <=32'hFFC00083;14'd11414:data <=32'hFFD60088;
14'd11415:data <=32'hFFED0088;14'd11416:data <=32'h00050083;14'd11417:data <=32'h001D0078;
14'd11418:data <=32'h00320065;14'd11419:data <=32'h0040004C;14'd11420:data <=32'h0045002F;
14'd11421:data <=32'h003E0013;14'd11422:data <=32'h002DFFFC;14'd11423:data <=32'h0016FFEE;
14'd11424:data <=32'hFFFCFFEC;14'd11425:data <=32'hFFE3FFF2;14'd11426:data <=32'hFFD10001;
14'd11427:data <=32'hFFC50015;14'd11428:data <=32'hFFC0002D;14'd11429:data <=32'hFFC40042;
14'd11430:data <=32'hFFCD0057;14'd11431:data <=32'hFFDA0069;14'd11432:data <=32'hFFEC0076;
14'd11433:data <=32'h00010080;14'd11434:data <=32'h001A0085;14'd11435:data <=32'h00320083;
14'd11436:data <=32'h004A007A;14'd11437:data <=32'h005F006B;14'd11438:data <=32'h006E0058;
14'd11439:data <=32'h00760043;14'd11440:data <=32'h0076002F;14'd11441:data <=32'h0071001F;
14'd11442:data <=32'h006B0016;14'd11443:data <=32'h00660014;14'd11444:data <=32'h00650014;
14'd11445:data <=32'h006B0014;14'd11446:data <=32'h00760011;14'd11447:data <=32'h00810009;
14'd11448:data <=32'h008EFFFA;14'd11449:data <=32'h0095FFE5;14'd11450:data <=32'h0098FFCE;
14'd11451:data <=32'h0095FFB7;14'd11452:data <=32'h008CFFA0;14'd11453:data <=32'h0081FF8B;
14'd11454:data <=32'h0073FF79;14'd11455:data <=32'h0061FF67;14'd11456:data <=32'h00D6FFCC;
14'd11457:data <=32'h00E4FF86;14'd11458:data <=32'h00CBFF4F;14'd11459:data <=32'h003DFF6C;
14'd11460:data <=32'hFFEEFF71;14'd11461:data <=32'hFFE0FF81;14'd11462:data <=32'hFFDAFF94;
14'd11463:data <=32'hFFDAFFA3;14'd11464:data <=32'hFFE2FFAC;14'd11465:data <=32'hFFEBFFAD;
14'd11466:data <=32'hFFF2FFA4;14'd11467:data <=32'hFFF1FF96;14'd11468:data <=32'hFFE6FF86;
14'd11469:data <=32'hFFD2FF7B;14'd11470:data <=32'hFFB8FF76;14'd11471:data <=32'hFF9CFF7A;
14'd11472:data <=32'hFF80FF88;14'd11473:data <=32'hFF69FF9C;14'd11474:data <=32'hFF57FFB6;
14'd11475:data <=32'hFF4AFFD3;14'd11476:data <=32'hFF42FFF3;14'd11477:data <=32'hFF440015;
14'd11478:data <=32'hFF4C0038;14'd11479:data <=32'hFF5D0059;14'd11480:data <=32'hFF770076;
14'd11481:data <=32'hFF9A008A;14'd11482:data <=32'hFFC10092;14'd11483:data <=32'hFFE7008E;
14'd11484:data <=32'h0009007D;14'd11485:data <=32'h00210064;14'd11486:data <=32'h002F0046;
14'd11487:data <=32'h00300029;14'd11488:data <=32'h00270011;14'd11489:data <=32'h001AFFFE;
14'd11490:data <=32'h0008FFF3;14'd11491:data <=32'hFFF7FFEE;14'd11492:data <=32'hFFE6FFEE;
14'd11493:data <=32'hFFD7FFF2;14'd11494:data <=32'hFFC8FFFA;14'd11495:data <=32'hFFBC0005;
14'd11496:data <=32'hFFB20013;14'd11497:data <=32'hFFAA0024;14'd11498:data <=32'hFFA70039;
14'd11499:data <=32'hFFA9004E;14'd11500:data <=32'hFFB10064;14'd11501:data <=32'hFFBE0077;
14'd11502:data <=32'hFFCE0086;14'd11503:data <=32'hFFE00092;14'd11504:data <=32'hFFF3009A;
14'd11505:data <=32'h000600A3;14'd11506:data <=32'h001C00A9;14'd11507:data <=32'h003300AF;
14'd11508:data <=32'h005000B2;14'd11509:data <=32'h007100AF;14'd11510:data <=32'h009600A4;
14'd11511:data <=32'h00BB008E;14'd11512:data <=32'h00D9006D;14'd11513:data <=32'h00F00043;
14'd11514:data <=32'h00F90013;14'd11515:data <=32'h00F7FFE4;14'd11516:data <=32'h00E8FFB7;
14'd11517:data <=32'h00D0FF93;14'd11518:data <=32'h00B2FF76;14'd11519:data <=32'h0093FF61;
14'd11520:data <=32'h009D0048;14'd11521:data <=32'h00CC0025;14'd11522:data <=32'h00E3FFE4;
14'd11523:data <=32'h0078FF5C;14'd11524:data <=32'h001AFF5E;14'd11525:data <=32'hFFFFFF72;
14'd11526:data <=32'hFFEFFF8D;14'd11527:data <=32'hFFE9FFA7;14'd11528:data <=32'hFFF0FFBE;
14'd11529:data <=32'hFFFFFFCC;14'd11530:data <=32'h0011FFD0;14'd11531:data <=32'h0022FFC6;
14'd11532:data <=32'h002AFFB6;14'd11533:data <=32'h0029FFA2;14'd11534:data <=32'h0020FF8E;
14'd11535:data <=32'h000FFF7F;14'd11536:data <=32'hFFF9FF76;14'd11537:data <=32'hFFE2FF73;
14'd11538:data <=32'hFFCCFF75;14'd11539:data <=32'hFFB4FF7B;14'd11540:data <=32'hFF9EFF86;
14'd11541:data <=32'hFF8AFF96;14'd11542:data <=32'hFF79FFAC;14'd11543:data <=32'hFF6EFFC7;
14'd11544:data <=32'hFF69FFE4;14'd11545:data <=32'hFF6D0002;14'd11546:data <=32'hFF7B001B;
14'd11547:data <=32'hFF8E002F;14'd11548:data <=32'hFFA3003A;14'd11549:data <=32'hFFB8003C;
14'd11550:data <=32'hFFCA003A;14'd11551:data <=32'hFFD60034;14'd11552:data <=32'hFFDE002E;
14'd11553:data <=32'hFFE30029;14'd11554:data <=32'hFFE90025;14'd11555:data <=32'hFFEE0022;
14'd11556:data <=32'hFFF3001C;14'd11557:data <=32'hFFF80014;14'd11558:data <=32'hFFFC0009;
14'd11559:data <=32'hFFFAFFFC;14'd11560:data <=32'hFFF3FFEF;14'd11561:data <=32'hFFE6FFE4;
14'd11562:data <=32'hFFD4FFDD;14'd11563:data <=32'hFFC0FFDD;14'd11564:data <=32'hFFA9FFE2;
14'd11565:data <=32'hFF96FFEF;14'd11566:data <=32'hFF830002;14'd11567:data <=32'hFF730018;
14'd11568:data <=32'hFF680035;14'd11569:data <=32'hFF610056;14'd11570:data <=32'hFF64007D;
14'd11571:data <=32'hFF6F00A6;14'd11572:data <=32'hFF8600D1;14'd11573:data <=32'hFFAC00F6;
14'd11574:data <=32'hFFDF0113;14'd11575:data <=32'h001A0121;14'd11576:data <=32'h0059011E;
14'd11577:data <=32'h00960109;14'd11578:data <=32'h00C900E4;14'd11579:data <=32'h00F100B4;
14'd11580:data <=32'h0109007E;14'd11581:data <=32'h01130047;14'd11582:data <=32'h01110014;
14'd11583:data <=32'h0105FFE4;14'd11584:data <=32'h008C0045;14'd11585:data <=32'h00AC0037;
14'd11586:data <=32'h00D5001E;14'd11587:data <=32'h0105FFD5;14'd11588:data <=32'h00B2FFB0;
14'd11589:data <=32'h0098FFA2;14'd11590:data <=32'h007FFF9C;14'd11591:data <=32'h006AFF9B;
14'd11592:data <=32'h005CFF9E;14'd11593:data <=32'h0054FFA1;14'd11594:data <=32'h0051FF9F;
14'd11595:data <=32'h004EFF98;14'd11596:data <=32'h0047FF8F;14'd11597:data <=32'h003BFF84;
14'd11598:data <=32'h002AFF7B;14'd11599:data <=32'h0015FF78;14'd11600:data <=32'h0000FF7B;
14'd11601:data <=32'hFFEFFF83;14'd11602:data <=32'hFFE0FF8F;14'd11603:data <=32'hFFD7FF9B;
14'd11604:data <=32'hFFD1FFA6;14'd11605:data <=32'hFFCDFFB0;14'd11606:data <=32'hFFCBFFB9;
14'd11607:data <=32'hFFC8FFC2;14'd11608:data <=32'hFFC8FFCC;14'd11609:data <=32'hFFCBFFD5;
14'd11610:data <=32'hFFCFFFDC;14'd11611:data <=32'hFFD4FFDF;14'd11612:data <=32'hFFD9FFDE;
14'd11613:data <=32'hFFDBFFDA;14'd11614:data <=32'hFFD9FFD3;14'd11615:data <=32'hFFD3FFD0;
14'd11616:data <=32'hFFC8FFD0;14'd11617:data <=32'hFFBCFFD4;14'd11618:data <=32'hFFB3FFE0;
14'd11619:data <=32'hFFAFFFEF;14'd11620:data <=32'hFFB1FFFF;14'd11621:data <=32'hFFBB000C;
14'd11622:data <=32'hFFC90014;14'd11623:data <=32'hFFD80015;14'd11624:data <=32'hFFE5000F;
14'd11625:data <=32'hFFEE0003;14'd11626:data <=32'hFFF1FFF5;14'd11627:data <=32'hFFEDFFE7;
14'd11628:data <=32'hFFE4FFDA;14'd11629:data <=32'hFFD6FFCE;14'd11630:data <=32'hFFC2FFC8;
14'd11631:data <=32'hFFADFFC6;14'd11632:data <=32'hFF93FFCA;14'd11633:data <=32'hFF79FFD6;
14'd11634:data <=32'hFF5FFFEC;14'd11635:data <=32'hFF49000A;14'd11636:data <=32'hFF3C0032;
14'd11637:data <=32'hFF3A0060;14'd11638:data <=32'hFF46008F;14'd11639:data <=32'hFF6100BB;
14'd11640:data <=32'hFF8600DD;14'd11641:data <=32'hFFB300F3;14'd11642:data <=32'hFFE300FD;
14'd11643:data <=32'h001000FA;14'd11644:data <=32'h003800EF;14'd11645:data <=32'h005A00DE;
14'd11646:data <=32'h007700C9;14'd11647:data <=32'h008F00B3;14'd11648:data <=32'h009B00B3;
14'd11649:data <=32'h00C100A0;14'd11650:data <=32'h00D80092;14'd11651:data <=32'h00AD00BB;
14'd11652:data <=32'h008A009D;14'd11653:data <=32'h009F008C;14'd11654:data <=32'h00B20078;
14'd11655:data <=32'h00C30061;14'd11656:data <=32'h00D30048;14'd11657:data <=32'h00E1002A;
14'd11658:data <=32'h00EC0007;14'd11659:data <=32'h00F0FFDE;14'd11660:data <=32'h00E8FFB1;
14'd11661:data <=32'h00D4FF86;14'd11662:data <=32'h00B3FF5F;14'd11663:data <=32'h0089FF46;
14'd11664:data <=32'h005AFF39;14'd11665:data <=32'h002CFF39;14'd11666:data <=32'h0003FF47;
14'd11667:data <=32'hFFE2FF5D;14'd11668:data <=32'hFFCDFF77;14'd11669:data <=32'hFFBEFF94;
14'd11670:data <=32'hFFB8FFB0;14'd11671:data <=32'hFFB8FFCA;14'd11672:data <=32'hFFBFFFE1;
14'd11673:data <=32'hFFCDFFF5;14'd11674:data <=32'hFFDF0002;14'd11675:data <=32'hFFF30009;
14'd11676:data <=32'h00090006;14'd11677:data <=32'h001CFFFB;14'd11678:data <=32'h0028FFE9;
14'd11679:data <=32'h002BFFD4;14'd11680:data <=32'h0026FFC0;14'd11681:data <=32'h0019FFB0;
14'd11682:data <=32'h0007FFA7;14'd11683:data <=32'hFFF4FFA6;14'd11684:data <=32'hFFE6FFAB;
14'd11685:data <=32'hFFDBFFB3;14'd11686:data <=32'hFFD5FFBB;14'd11687:data <=32'hFFD3FFC1;
14'd11688:data <=32'hFFD2FFC5;14'd11689:data <=32'hFFD2FFC6;14'd11690:data <=32'hFFCFFFC6;
14'd11691:data <=32'hFFCAFFC5;14'd11692:data <=32'hFFC3FFC5;14'd11693:data <=32'hFFBBFFC7;
14'd11694:data <=32'hFFB5FFC9;14'd11695:data <=32'hFFADFFCC;14'd11696:data <=32'hFFA3FFD0;
14'd11697:data <=32'hFF99FFD5;14'd11698:data <=32'hFF8EFFDC;14'd11699:data <=32'hFF81FFE7;
14'd11700:data <=32'hFF76FFF7;14'd11701:data <=32'hFF6F000C;14'd11702:data <=32'hFF6D0024;
14'd11703:data <=32'hFF72003C;14'd11704:data <=32'hFF7D004F;14'd11705:data <=32'hFF8D005E;
14'd11706:data <=32'hFF9C0066;14'd11707:data <=32'hFFA8006A;14'd11708:data <=32'hFFB0006D;
14'd11709:data <=32'hFFB20070;14'd11710:data <=32'hFFB40078;14'd11711:data <=32'hFFB80086;
14'd11712:data <=32'hFFE30103;14'd11713:data <=32'h00120113;14'd11714:data <=32'h00320103;
14'd11715:data <=32'hFFD100B4;14'd11716:data <=32'hFFAC00BE;14'd11717:data <=32'hFFC800D8;
14'd11718:data <=32'hFFEB00EC;14'd11719:data <=32'h001400F9;14'd11720:data <=32'h004300FE;
14'd11721:data <=32'h007600F7;14'd11722:data <=32'h00AA00E4;14'd11723:data <=32'h00DA00C1;
14'd11724:data <=32'h00FF0090;14'd11725:data <=32'h01170056;14'd11726:data <=32'h011D0018;
14'd11727:data <=32'h010FFFDC;14'd11728:data <=32'h00F3FFA9;14'd11729:data <=32'h00CDFF81;
14'd11730:data <=32'h00A2FF69;14'd11731:data <=32'h0077FF5C;14'd11732:data <=32'h004FFF5B;
14'd11733:data <=32'h0029FF61;14'd11734:data <=32'h000BFF6F;14'd11735:data <=32'hFFF1FF81;
14'd11736:data <=32'hFFDDFF98;14'd11737:data <=32'hFFD0FFB2;14'd11738:data <=32'hFFCCFFCD;
14'd11739:data <=32'hFFD1FFE7;14'd11740:data <=32'hFFDDFFFC;14'd11741:data <=32'hFFEE0009;
14'd11742:data <=32'h0003000F;14'd11743:data <=32'h0016000E;14'd11744:data <=32'h00240007;
14'd11745:data <=32'h002DFFFD;14'd11746:data <=32'h0033FFF2;14'd11747:data <=32'h0037FFE9;
14'd11748:data <=32'h003AFFE1;14'd11749:data <=32'h003DFFD9;14'd11750:data <=32'h0042FFCC;
14'd11751:data <=32'h0045FFBE;14'd11752:data <=32'h0044FFAB;14'd11753:data <=32'h003DFF96;
14'd11754:data <=32'h0031FF81;14'd11755:data <=32'h001CFF6F;14'd11756:data <=32'h0002FF62;
14'd11757:data <=32'hFFE4FF5D;14'd11758:data <=32'hFFC6FF60;14'd11759:data <=32'hFFA9FF6A;
14'd11760:data <=32'hFF90FF79;14'd11761:data <=32'hFF7CFF8D;14'd11762:data <=32'hFF6CFFA4;
14'd11763:data <=32'hFF60FFBD;14'd11764:data <=32'hFF5AFFD9;14'd11765:data <=32'hFF5AFFF6;
14'd11766:data <=32'hFF610012;14'd11767:data <=32'hFF71002B;14'd11768:data <=32'hFF85003B;
14'd11769:data <=32'hFF9E0043;14'd11770:data <=32'hFFB50040;14'd11771:data <=32'hFFC60035;
14'd11772:data <=32'hFFCD0025;14'd11773:data <=32'hFFC80014;14'd11774:data <=32'hFFBA000A;
14'd11775:data <=32'hFFA60008;14'd11776:data <=32'hFF5C005D;14'd11777:data <=32'hFF5D0080;
14'd11778:data <=32'hFF790094;14'd11779:data <=32'hFFA90045;14'd11780:data <=32'hFF6C004B;
14'd11781:data <=32'hFF6D0069;14'd11782:data <=32'hFF760088;14'd11783:data <=32'hFF8700A5;
14'd11784:data <=32'hFF9F00C1;14'd11785:data <=32'hFFC000DA;14'd11786:data <=32'hFFEA00E9;
14'd11787:data <=32'h001800EE;14'd11788:data <=32'h004700E5;14'd11789:data <=32'h007100CF;
14'd11790:data <=32'h009200AF;14'd11791:data <=32'h00A70089;14'd11792:data <=32'h00B10063;
14'd11793:data <=32'h00B00041;14'd11794:data <=32'h00AB0023;14'd11795:data <=32'h00A1000C;
14'd11796:data <=32'h0097FFF8;14'd11797:data <=32'h008CFFE6;14'd11798:data <=32'h0081FFD7;
14'd11799:data <=32'h0072FFC9;14'd11800:data <=32'h0061FFBC;14'd11801:data <=32'h004EFFB7;
14'd11802:data <=32'h003BFFB5;14'd11803:data <=32'h0028FFB6;14'd11804:data <=32'h001AFFBE;
14'd11805:data <=32'h000EFFC7;14'd11806:data <=32'h0006FFD1;14'd11807:data <=32'h0001FFDA;
14'd11808:data <=32'hFFFCFFE4;14'd11809:data <=32'hFFFAFFF0;14'd11810:data <=32'hFFF9FFFD;
14'd11811:data <=32'hFFFE000B;14'd11812:data <=32'h0008001B;14'd11813:data <=32'h001A0029;
14'd11814:data <=32'h0031002F;14'd11815:data <=32'h004F002D;14'd11816:data <=32'h006B0020;
14'd11817:data <=32'h00840007;14'd11818:data <=32'h0094FFE7;14'd11819:data <=32'h009AFFC0;
14'd11820:data <=32'h0094FF98;14'd11821:data <=32'h0082FF73;14'd11822:data <=32'h0068FF55;
14'd11823:data <=32'h0047FF3F;14'd11824:data <=32'h0021FF31;14'd11825:data <=32'hFFFBFF2D;
14'd11826:data <=32'hFFD5FF2F;14'd11827:data <=32'hFFB1FF3C;14'd11828:data <=32'hFF8FFF4E;
14'd11829:data <=32'hFF74FF69;14'd11830:data <=32'hFF61FF89;14'd11831:data <=32'hFF58FFAC;
14'd11832:data <=32'hFF59FFCE;14'd11833:data <=32'hFF64FFE9;14'd11834:data <=32'hFF75FFFD;
14'd11835:data <=32'hFF880006;14'd11836:data <=32'hFF960007;14'd11837:data <=32'hFF9D0002;
14'd11838:data <=32'hFF9DFFFC;14'd11839:data <=32'hFF95FFF9;14'd11840:data <=32'hFFB5FFE0;
14'd11841:data <=32'hFF9BFFDC;14'd11842:data <=32'hFF89FFF1;14'd11843:data <=32'hFF86003F;
14'd11844:data <=32'hFF550041;14'd11845:data <=32'hFF620058;14'd11846:data <=32'hFF71006D;
14'd11847:data <=32'hFF84007D;14'd11848:data <=32'hFF98008A;14'd11849:data <=32'hFFAD0096;
14'd11850:data <=32'hFFC5009D;14'd11851:data <=32'hFFDF009E;14'd11852:data <=32'hFFF9009A;
14'd11853:data <=32'h0010008E;14'd11854:data <=32'h0020007D;14'd11855:data <=32'h0029006A;
14'd11856:data <=32'h002A005A;14'd11857:data <=32'h0025004F;14'd11858:data <=32'h001F004C;
14'd11859:data <=32'h001C004E;14'd11860:data <=32'h001E0055;14'd11861:data <=32'h0027005B;
14'd11862:data <=32'h0034005D;14'd11863:data <=32'h0043005A;14'd11864:data <=32'h00520051;
14'd11865:data <=32'h005F0043;14'd11866:data <=32'h00660033;14'd11867:data <=32'h006B0022;
14'd11868:data <=32'h006B0010;14'd11869:data <=32'h0067FFFF;14'd11870:data <=32'h0060FFEF;
14'd11871:data <=32'h0055FFE1;14'd11872:data <=32'h0045FFD5;14'd11873:data <=32'h0031FFCE;
14'd11874:data <=32'h001DFFD0;14'd11875:data <=32'h0008FFD9;14'd11876:data <=32'hFFF9FFEA;
14'd11877:data <=32'hFFF20001;14'd11878:data <=32'hFFF5001A;14'd11879:data <=32'h00030031;
14'd11880:data <=32'h00190042;14'd11881:data <=32'h00350048;14'd11882:data <=32'h00530044;
14'd11883:data <=32'h006D0036;14'd11884:data <=32'h00820021;14'd11885:data <=32'h00910009;
14'd11886:data <=32'h0098FFEC;14'd11887:data <=32'h0099FFD2;14'd11888:data <=32'h0095FFB8;
14'd11889:data <=32'h008DFF9D;14'd11890:data <=32'h0081FF85;14'd11891:data <=32'h0070FF6F;
14'd11892:data <=32'h005AFF5B;14'd11893:data <=32'h0041FF4D;14'd11894:data <=32'h0025FF45;
14'd11895:data <=32'h000AFF42;14'd11896:data <=32'hFFF1FF44;14'd11897:data <=32'hFFDCFF49;
14'd11898:data <=32'hFFC9FF4E;14'd11899:data <=32'hFFB8FF53;14'd11900:data <=32'hFFA4FF56;
14'd11901:data <=32'hFF8DFF5B;14'd11902:data <=32'hFF73FF63;14'd11903:data <=32'hFF55FF73;
14'd11904:data <=32'hFFDAFFEF;14'd11905:data <=32'hFFD6FFD8;14'd11906:data <=32'hFFBAFFC2;
14'd11907:data <=32'hFF27FFBA;14'd11908:data <=32'hFEE9FFD8;14'd11909:data <=32'hFEEE000E;
14'd11910:data <=32'hFF00003F;14'd11911:data <=32'hFF1D0067;14'd11912:data <=32'hFF3E0087;
14'd11913:data <=32'hFF63009E;14'd11914:data <=32'hFF8C00AC;14'd11915:data <=32'hFFB500AF;
14'd11916:data <=32'hFFDD00A9;14'd11917:data <=32'h00010096;14'd11918:data <=32'h0018007C;
14'd11919:data <=32'h0026005D;14'd11920:data <=32'h0025003E;14'd11921:data <=32'h001A0027;
14'd11922:data <=32'h00080019;14'd11923:data <=32'hFFF30016;14'd11924:data <=32'hFFE2001D;
14'd11925:data <=32'hFFD9002B;14'd11926:data <=32'hFFD6003B;14'd11927:data <=32'hFFDC004B;
14'd11928:data <=32'hFFE60057;14'd11929:data <=32'hFFF30060;14'd11930:data <=32'h00010064;
14'd11931:data <=32'h00100064;14'd11932:data <=32'h001E0062;14'd11933:data <=32'h002D005C;
14'd11934:data <=32'h003A0053;14'd11935:data <=32'h00450047;14'd11936:data <=32'h004C0038;
14'd11937:data <=32'h004D0027;14'd11938:data <=32'h00490017;14'd11939:data <=32'h0040000C;
14'd11940:data <=32'h00330007;14'd11941:data <=32'h00280007;14'd11942:data <=32'h0020000E;
14'd11943:data <=32'h001C0016;14'd11944:data <=32'h001E001F;14'd11945:data <=32'h00240026;
14'd11946:data <=32'h002C0027;14'd11947:data <=32'h00340026;14'd11948:data <=32'h003B0023;
14'd11949:data <=32'h003E0020;14'd11950:data <=32'h0042001F;14'd11951:data <=32'h0045001F;
14'd11952:data <=32'h004A0020;14'd11953:data <=32'h00540023;14'd11954:data <=32'h00620022;
14'd11955:data <=32'h0072001D;14'd11956:data <=32'h00840010;14'd11957:data <=32'h00940001;
14'd11958:data <=32'h00A0FFEA;14'd11959:data <=32'h00A9FFD1;14'd11960:data <=32'h00AFFFB4;
14'd11961:data <=32'h00B0FF94;14'd11962:data <=32'h00ABFF70;14'd11963:data <=32'h009EFF4B;
14'd11964:data <=32'h0088FF23;14'd11965:data <=32'h0065FEFD;14'd11966:data <=32'h0035FEDE;
14'd11967:data <=32'hFFFBFECC;14'd11968:data <=32'hFFDFFF98;14'd11969:data <=32'hFFD7FF87;
14'd11970:data <=32'hFFD6FF6A;14'd11971:data <=32'hFFAEFEF5;14'd11972:data <=32'hFF44FF00;
14'd11973:data <=32'hFF1DFF30;14'd11974:data <=32'hFF04FF65;14'd11975:data <=32'hFEF9FF9B;
14'd11976:data <=32'hFEF8FFCE;14'd11977:data <=32'hFF02FFFF;14'd11978:data <=32'hFF15002B;
14'd11979:data <=32'hFF300050;14'd11980:data <=32'hFF53006B;14'd11981:data <=32'hFF79007B;
14'd11982:data <=32'hFF9F007E;14'd11983:data <=32'hFFC00076;14'd11984:data <=32'hFFD80068;
14'd11985:data <=32'hFFE60055;14'd11986:data <=32'hFFEA0045;14'd11987:data <=32'hFFE9003A;
14'd11988:data <=32'hFFE60034;14'd11989:data <=32'hFFE40033;14'd11990:data <=32'hFFE40034;
14'd11991:data <=32'hFFE70035;14'd11992:data <=32'hFFEB0034;14'd11993:data <=32'hFFEE0032;
14'd11994:data <=32'hFFEF002E;14'd11995:data <=32'hFFEE002B;14'd11996:data <=32'hFFEB002B;
14'd11997:data <=32'hFFE7002D;14'd11998:data <=32'hFFE60031;14'd11999:data <=32'hFFE60038;
14'd12000:data <=32'hFFE9003D;14'd12001:data <=32'hFFEC0040;14'd12002:data <=32'hFFF10043;
14'd12003:data <=32'hFFF40048;14'd12004:data <=32'hFFF8004D;14'd12005:data <=32'hFFFE0053;
14'd12006:data <=32'h00060059;14'd12007:data <=32'h0013005F;14'd12008:data <=32'h0022005F;
14'd12009:data <=32'h0033005C;14'd12010:data <=32'h00420051;14'd12011:data <=32'h004D0042;
14'd12012:data <=32'h00510030;14'd12013:data <=32'h004E001E;14'd12014:data <=32'h00440011;
14'd12015:data <=32'h0036000C;14'd12016:data <=32'h0028000E;14'd12017:data <=32'h001D0018;
14'd12018:data <=32'h001A0027;14'd12019:data <=32'h001E0037;14'd12020:data <=32'h002B0047;
14'd12021:data <=32'h003D0052;14'd12022:data <=32'h00530058;14'd12023:data <=32'h006F0057;
14'd12024:data <=32'h008D0050;14'd12025:data <=32'h00AA0041;14'd12026:data <=32'h00C70028;
14'd12027:data <=32'h00E10004;14'd12028:data <=32'h00F3FFD7;14'd12029:data <=32'h00F9FFA2;
14'd12030:data <=32'h00EEFF69;14'd12031:data <=32'h00D3FF32;14'd12032:data <=32'h0096FF77;
14'd12033:data <=32'h008CFF48;14'd12034:data <=32'h0084FF2D;14'd12035:data <=32'h008DFF33;
14'd12036:data <=32'h002FFF11;14'd12037:data <=32'h0007FF15;14'd12038:data <=32'hFFE6FF1E;
14'd12039:data <=32'hFFCAFF2C;14'd12040:data <=32'hFFB0FF3B;14'd12041:data <=32'hFF98FF4C;
14'd12042:data <=32'hFF84FF61;14'd12043:data <=32'hFF73FF79;14'd12044:data <=32'hFF68FF93;
14'd12045:data <=32'hFF62FFAB;14'd12046:data <=32'hFF62FFC2;14'd12047:data <=32'hFF64FFD7;
14'd12048:data <=32'hFF67FFE7;14'd12049:data <=32'hFF69FFF6;14'd12050:data <=32'hFF6A0007;
14'd12051:data <=32'hFF6C001B;14'd12052:data <=32'hFF720031;14'd12053:data <=32'hFF7F0047;
14'd12054:data <=32'hFF93005B;14'd12055:data <=32'hFFAC0068;14'd12056:data <=32'hFFCB006C;
14'd12057:data <=32'hFFE60066;14'd12058:data <=32'hFFFE0058;14'd12059:data <=32'h000D0044;
14'd12060:data <=32'h0013002E;14'd12061:data <=32'h00120019;14'd12062:data <=32'h000B0008;
14'd12063:data <=32'hFFFFFFFB;14'd12064:data <=32'hFFF1FFF3;14'd12065:data <=32'hFFE1FFF1;
14'd12066:data <=32'hFFCFFFF2;14'd12067:data <=32'hFFBEFFFA;14'd12068:data <=32'hFFB00007;
14'd12069:data <=32'hFFA5001A;14'd12070:data <=32'hFFA00032;14'd12071:data <=32'hFFA3004B;
14'd12072:data <=32'hFFAF0063;14'd12073:data <=32'hFFC20076;14'd12074:data <=32'hFFDC0082;
14'd12075:data <=32'hFFF50084;14'd12076:data <=32'h000D007E;14'd12077:data <=32'h001F0072;
14'd12078:data <=32'h00290065;14'd12079:data <=32'h002C0057;14'd12080:data <=32'h002A004F;
14'd12081:data <=32'h0028004C;14'd12082:data <=32'h0026004D;14'd12083:data <=32'h00280052;
14'd12084:data <=32'h002E0057;14'd12085:data <=32'h0038005C;14'd12086:data <=32'h0044005F;
14'd12087:data <=32'h0051005F;14'd12088:data <=32'h0061005D;14'd12089:data <=32'h00730059;
14'd12090:data <=32'h00870052;14'd12091:data <=32'h009B0044;14'd12092:data <=32'h00B10030;
14'd12093:data <=32'h00C00014;14'd12094:data <=32'h00C9FFF2;14'd12095:data <=32'h00C8FFCD;
14'd12096:data <=32'h00F5003B;14'd12097:data <=32'h011C0002;14'd12098:data <=32'h011AFFCC;
14'd12099:data <=32'h0099FFC1;14'd12100:data <=32'h0056FFA3;14'd12101:data <=32'h004DFFA7;
14'd12102:data <=32'h004AFFAB;14'd12103:data <=32'h004CFFAC;14'd12104:data <=32'h004FFFA4;
14'd12105:data <=32'h0050FF98;14'd12106:data <=32'h004BFF88;14'd12107:data <=32'h0043FF77;
14'd12108:data <=32'h0034FF69;14'd12109:data <=32'h0021FF5B;14'd12110:data <=32'h000CFF50;
14'd12111:data <=32'hFFF3FF48;14'd12112:data <=32'hFFD6FF45;14'd12113:data <=32'hFFB5FF46;
14'd12114:data <=32'hFF91FF51;14'd12115:data <=32'hFF6EFF66;14'd12116:data <=32'hFF52FF87;
14'd12117:data <=32'hFF3EFFAF;14'd12118:data <=32'hFF38FFDD;14'd12119:data <=32'hFF41000A;
14'd12120:data <=32'hFF550030;14'd12121:data <=32'hFF74004D;14'd12122:data <=32'hFF97005D;
14'd12123:data <=32'hFFB90061;14'd12124:data <=32'hFFD9005C;14'd12125:data <=32'hFFF10050;
14'd12126:data <=32'h0003003E;14'd12127:data <=32'h0010002B;14'd12128:data <=32'h00150016;
14'd12129:data <=32'h00150001;14'd12130:data <=32'h000FFFED;14'd12131:data <=32'h0002FFDC;
14'd12132:data <=32'hFFF0FFD0;14'd12133:data <=32'hFFDAFFCA;14'd12134:data <=32'hFFC2FFCC;
14'd12135:data <=32'hFFACFFD5;14'd12136:data <=32'hFF9BFFE5;14'd12137:data <=32'hFF90FFF9;
14'd12138:data <=32'hFF8A000E;14'd12139:data <=32'hFF8A0021;14'd12140:data <=32'hFF8E0031;
14'd12141:data <=32'hFF910040;14'd12142:data <=32'hFF94004F;14'd12143:data <=32'hFF98005D;
14'd12144:data <=32'hFF9C0070;14'd12145:data <=32'hFFA30085;14'd12146:data <=32'hFFB1009C;
14'd12147:data <=32'hFFC600B0;14'd12148:data <=32'hFFE200C2;14'd12149:data <=32'h000300CC;
14'd12150:data <=32'h002800CE;14'd12151:data <=32'h004B00C7;14'd12152:data <=32'h006B00B9;
14'd12153:data <=32'h008700A4;14'd12154:data <=32'h009F008C;14'd12155:data <=32'h00B20070;
14'd12156:data <=32'h00C00051;14'd12157:data <=32'h00C7002F;14'd12158:data <=32'h00C7000B;
14'd12159:data <=32'h00BDFFE8;14'd12160:data <=32'h007300B1;14'd12161:data <=32'h00AD00A4;
14'd12162:data <=32'h00DA0074;14'd12163:data <=32'h009DFFD4;14'd12164:data <=32'h004FFFB7;
14'd12165:data <=32'h003BFFC6;14'd12166:data <=32'h0032FFD9;14'd12167:data <=32'h0034FFEA;
14'd12168:data <=32'h0040FFF5;14'd12169:data <=32'h004EFFF8;14'd12170:data <=32'h005DFFF3;
14'd12171:data <=32'h006AFFE7;14'd12172:data <=32'h0073FFD7;14'd12173:data <=32'h0078FFC3;
14'd12174:data <=32'h0079FFAC;14'd12175:data <=32'h0074FF93;14'd12176:data <=32'h0068FF79;
14'd12177:data <=32'h0053FF60;14'd12178:data <=32'h0036FF4B;14'd12179:data <=32'h0012FF3F;
14'd12180:data <=32'hFFEAFF3E;14'd12181:data <=32'hFFC4FF4A;14'd12182:data <=32'hFFA3FF61;
14'd12183:data <=32'hFF8CFF7F;14'd12184:data <=32'hFF80FF9F;14'd12185:data <=32'hFF7EFFBF;
14'd12186:data <=32'hFF83FFDB;14'd12187:data <=32'hFF8EFFF0;14'd12188:data <=32'hFF9AFFFF;
14'd12189:data <=32'hFFA7000A;14'd12190:data <=32'hFFB40014;14'd12191:data <=32'hFFC10019;
14'd12192:data <=32'hFFCF001D;14'd12193:data <=32'hFFDF001E;14'd12194:data <=32'hFFEC001A;
14'd12195:data <=32'hFFF90013;14'd12196:data <=32'h00030006;14'd12197:data <=32'h0007FFF7;
14'd12198:data <=32'h0007FFE7;14'd12199:data <=32'h0002FFD9;14'd12200:data <=32'hFFFAFFCD;
14'd12201:data <=32'hFFEEFFC3;14'd12202:data <=32'hFFE0FFB9;14'd12203:data <=32'hFFD1FFB2;
14'd12204:data <=32'hFFBFFFAD;14'd12205:data <=32'hFFA6FFAB;14'd12206:data <=32'hFF8AFFAE;
14'd12207:data <=32'hFF6BFFBA;14'd12208:data <=32'hFF4CFFD0;14'd12209:data <=32'hFF30FFF1;
14'd12210:data <=32'hFF1E001E;14'd12211:data <=32'hFF190051;14'd12212:data <=32'hFF220086;
14'd12213:data <=32'hFF3B00B8;14'd12214:data <=32'hFF5F00E2;14'd12215:data <=32'hFF8F0101;
14'd12216:data <=32'hFFC20113;14'd12217:data <=32'hFFF70119;14'd12218:data <=32'h002B0114;
14'd12219:data <=32'h005D0104;14'd12220:data <=32'h008900E9;14'd12221:data <=32'h00AE00C6;
14'd12222:data <=32'h00C9009A;14'd12223:data <=32'h00D7006A;14'd12224:data <=32'h003B0090;
14'd12225:data <=32'h005A0094;14'd12226:data <=32'h00880091;14'd12227:data <=32'h00D20055;
14'd12228:data <=32'h0093001D;14'd12229:data <=32'h00850013;14'd12230:data <=32'h007B000D;
14'd12231:data <=32'h0076000D;14'd12232:data <=32'h0077000A;14'd12233:data <=32'h007A0004;
14'd12234:data <=32'h007DFFF9;14'd12235:data <=32'h007CFFED;14'd12236:data <=32'h007BFFE0;
14'd12237:data <=32'h0076FFD4;14'd12238:data <=32'h0071FFC8;14'd12239:data <=32'h006AFFBE;
14'd12240:data <=32'h0063FFB2;14'd12241:data <=32'h005BFFA7;14'd12242:data <=32'h004FFF9B;
14'd12243:data <=32'h003EFF92;14'd12244:data <=32'h002BFF8E;14'd12245:data <=32'h0017FF8F;
14'd12246:data <=32'h0007FF96;14'd12247:data <=32'hFFFAFFA2;14'd12248:data <=32'hFFF4FFAE;
14'd12249:data <=32'hFFF3FFB7;14'd12250:data <=32'hFFF6FFBD;14'd12251:data <=32'hFFF9FFBE;
14'd12252:data <=32'hFFF8FFBB;14'd12253:data <=32'hFFF3FFB7;14'd12254:data <=32'hFFEBFFB4;
14'd12255:data <=32'hFFE0FFB7;14'd12256:data <=32'hFFD5FFBD;14'd12257:data <=32'hFFCDFFC7;
14'd12258:data <=32'hFFC9FFD3;14'd12259:data <=32'hFFCCFFE0;14'd12260:data <=32'hFFD0FFEA;
14'd12261:data <=32'hFFD8FFF3;14'd12262:data <=32'hFFE2FFF7;14'd12263:data <=32'hFFECFFF8;
14'd12264:data <=32'hFFF6FFF6;14'd12265:data <=32'h0000FFF0;14'd12266:data <=32'h000BFFE5;
14'd12267:data <=32'h0012FFD5;14'd12268:data <=32'h0013FFC0;14'd12269:data <=32'h000CFFA8;
14'd12270:data <=32'hFFFDFF8F;14'd12271:data <=32'hFFE0FF7A;14'd12272:data <=32'hFFBCFF6E;
14'd12273:data <=32'hFF91FF6D;14'd12274:data <=32'hFF66FF7C;14'd12275:data <=32'hFF3EFF98;
14'd12276:data <=32'hFF20FFBF;14'd12277:data <=32'hFF0EFFED;14'd12278:data <=32'hFF09001E;
14'd12279:data <=32'hFF0F004D;14'd12280:data <=32'hFF200078;14'd12281:data <=32'hFF38009E;
14'd12282:data <=32'hFF5600BD;14'd12283:data <=32'hFF7900D7;14'd12284:data <=32'hFFA000E9;
14'd12285:data <=32'hFFC900F2;14'd12286:data <=32'hFFF300F2;14'd12287:data <=32'h001B00E8;
14'd12288:data <=32'h002500CF;14'd12289:data <=32'h004500CD;14'd12290:data <=32'h005700CE;
14'd12291:data <=32'h002B00EF;14'd12292:data <=32'h001200CB;14'd12293:data <=32'h002900CD;
14'd12294:data <=32'h004500CD;14'd12295:data <=32'h006500CA;14'd12296:data <=32'h008800BC;
14'd12297:data <=32'h00AA00A4;14'd12298:data <=32'h00C60083;14'd12299:data <=32'h00D9005A;
14'd12300:data <=32'h00E0002F;14'd12301:data <=32'h00DB0004;14'd12302:data <=32'h00CEFFDF;
14'd12303:data <=32'h00B9FFBF;14'd12304:data <=32'h00A0FFA7;14'd12305:data <=32'h0084FF95;
14'd12306:data <=32'h0066FF89;14'd12307:data <=32'h0047FF84;14'd12308:data <=32'h0028FF88;
14'd12309:data <=32'h000CFF94;14'd12310:data <=32'hFFF7FFA8;14'd12311:data <=32'hFFEBFFC1;
14'd12312:data <=32'hFFE9FFDB;14'd12313:data <=32'hFFF2FFF1;14'd12314:data <=32'h00020000;
14'd12315:data <=32'h00160007;14'd12316:data <=32'h002A0002;14'd12317:data <=32'h0038FFF6;
14'd12318:data <=32'h003FFFE6;14'd12319:data <=32'h003FFFD5;14'd12320:data <=32'h0039FFC7;
14'd12321:data <=32'h0030FFBD;14'd12322:data <=32'h0025FFB7;14'd12323:data <=32'h001BFFB5;
14'd12324:data <=32'h0012FFB4;14'd12325:data <=32'h0009FFB5;14'd12326:data <=32'h0003FFB8;
14'd12327:data <=32'hFFFDFFBB;14'd12328:data <=32'hFFFAFFBF;14'd12329:data <=32'hFFF7FFC3;
14'd12330:data <=32'hFFF8FFC7;14'd12331:data <=32'hFFFCFFC7;14'd12332:data <=32'h0002FFC5;
14'd12333:data <=32'h0005FFBD;14'd12334:data <=32'h0005FFB0;14'd12335:data <=32'hFFFFFFA1;
14'd12336:data <=32'hFFF1FF93;14'd12337:data <=32'hFFDDFF87;14'd12338:data <=32'hFFC5FF84;
14'd12339:data <=32'hFFACFF89;14'd12340:data <=32'hFF95FF95;14'd12341:data <=32'hFF84FFA6;
14'd12342:data <=32'hFF78FFB9;14'd12343:data <=32'hFF71FFCA;14'd12344:data <=32'hFF6EFFDA;
14'd12345:data <=32'hFF69FFE8;14'd12346:data <=32'hFF64FFF6;14'd12347:data <=32'hFF5F0004;
14'd12348:data <=32'hFF5B0015;14'd12349:data <=32'hFF570029;14'd12350:data <=32'hFF580040;
14'd12351:data <=32'hFF5C0055;14'd12352:data <=32'hFF7500CE;14'd12353:data <=32'hFF9600E4;
14'd12354:data <=32'hFFAF00DD;14'd12355:data <=32'hFF5F007A;14'd12356:data <=32'hFF32007C;
14'd12357:data <=32'hFF3D00A9;14'd12358:data <=32'hFF5600D6;14'd12359:data <=32'hFF7B00FF;
14'd12360:data <=32'hFFAE011F;14'd12361:data <=32'hFFEB012F;14'd12362:data <=32'h002C012D;
14'd12363:data <=32'h00690119;14'd12364:data <=32'h009B00F6;14'd12365:data <=32'h00C200CB;
14'd12366:data <=32'h00DB009A;14'd12367:data <=32'h00E70066;14'd12368:data <=32'h00E90035;
14'd12369:data <=32'h00DF0007;14'd12370:data <=32'h00CDFFDE;14'd12371:data <=32'h00B2FFBC;
14'd12372:data <=32'h008FFFA1;14'd12373:data <=32'h0069FF92;14'd12374:data <=32'h0041FF91;
14'd12375:data <=32'h001FFF9B;14'd12376:data <=32'h0004FFAF;14'd12377:data <=32'hFFF4FFC7;
14'd12378:data <=32'hFFEFFFE1;14'd12379:data <=32'hFFF3FFF7;14'd12380:data <=32'hFFFD0007;
14'd12381:data <=32'h00090010;14'd12382:data <=32'h00160013;14'd12383:data <=32'h00200014;
14'd12384:data <=32'h00280013;14'd12385:data <=32'h002F0011;14'd12386:data <=32'h0038000F;
14'd12387:data <=32'h0041000C;14'd12388:data <=32'h004C0006;14'd12389:data <=32'h0056FFFD;
14'd12390:data <=32'h005EFFEF;14'd12391:data <=32'h0063FFDF;14'd12392:data <=32'h0064FFCE;
14'd12393:data <=32'h0061FFBC;14'd12394:data <=32'h005AFFAB;14'd12395:data <=32'h0051FF9D;
14'd12396:data <=32'h0046FF90;14'd12397:data <=32'h0039FF83;14'd12398:data <=32'h0029FF77;
14'd12399:data <=32'h0016FF6E;14'd12400:data <=32'hFFFDFF68;14'd12401:data <=32'hFFE4FF67;
14'd12402:data <=32'hFFCAFF6E;14'd12403:data <=32'hFFB2FF7D;14'd12404:data <=32'hFFA1FF93;
14'd12405:data <=32'hFF99FFAC;14'd12406:data <=32'hFF9AFFC3;14'd12407:data <=32'hFFA3FFD5;
14'd12408:data <=32'hFFB0FFDF;14'd12409:data <=32'hFFBEFFE0;14'd12410:data <=32'hFFC6FFDA;
14'd12411:data <=32'hFFC9FFCF;14'd12412:data <=32'hFFC3FFC3;14'd12413:data <=32'hFFB8FFB9;
14'd12414:data <=32'hFFA7FFB2;14'd12415:data <=32'hFF94FFB1;14'd12416:data <=32'hFF3EFFFB;
14'd12417:data <=32'hFF330015;14'd12418:data <=32'hFF440025;14'd12419:data <=32'hFF7EFFDA;
14'd12420:data <=32'hFF35FFC9;14'd12421:data <=32'hFF1DFFEE;14'd12422:data <=32'hFF0F001C;
14'd12423:data <=32'hFF0D004F;14'd12424:data <=32'hFF1B0083;14'd12425:data <=32'hFF3A00B1;
14'd12426:data <=32'hFF6200D4;14'd12427:data <=32'hFF9200EA;14'd12428:data <=32'hFFC200F3;
14'd12429:data <=32'hFFEF00F0;14'd12430:data <=32'h001600E4;14'd12431:data <=32'h003800D2;
14'd12432:data <=32'h005500BD;14'd12433:data <=32'h006D00A5;14'd12434:data <=32'h007F0088;
14'd12435:data <=32'h008C006A;14'd12436:data <=32'h0090004B;14'd12437:data <=32'h008D002D;
14'd12438:data <=32'h00810013;14'd12439:data <=32'h0073FFFF;14'd12440:data <=32'h0062FFF4;
14'd12441:data <=32'h0053FFED;14'd12442:data <=32'h0046FFEA;14'd12443:data <=32'h003BFFE8;
14'd12444:data <=32'h0032FFE6;14'd12445:data <=32'h0029FFE5;14'd12446:data <=32'h001EFFE4;
14'd12447:data <=32'h0011FFE7;14'd12448:data <=32'h0004FFED;14'd12449:data <=32'hFFF8FFFB;
14'd12450:data <=32'hFFF2000D;14'd12451:data <=32'hFFF30023;14'd12452:data <=32'hFFFE0038;
14'd12453:data <=32'h00110049;14'd12454:data <=32'h00290053;14'd12455:data <=32'h00450055;
14'd12456:data <=32'h0061004E;14'd12457:data <=32'h007A0040;14'd12458:data <=32'h0090002A;
14'd12459:data <=32'h00A10011;14'd12460:data <=32'h00ACFFF2;14'd12461:data <=32'h00AFFFD1;
14'd12462:data <=32'h00ABFFAD;14'd12463:data <=32'h009FFF8A;14'd12464:data <=32'h0088FF6A;
14'd12465:data <=32'h0069FF50;14'd12466:data <=32'h0043FF40;14'd12467:data <=32'h001BFF3D;
14'd12468:data <=32'hFFF4FF44;14'd12469:data <=32'hFFD6FF57;14'd12470:data <=32'hFFC2FF70;
14'd12471:data <=32'hFFB8FF8A;14'd12472:data <=32'hFFB7FF9F;14'd12473:data <=32'hFFBEFFAE;
14'd12474:data <=32'hFFC6FFB7;14'd12475:data <=32'hFFCDFFB8;14'd12476:data <=32'hFFCFFFB4;
14'd12477:data <=32'hFFCFFFAF;14'd12478:data <=32'hFFC9FFA8;14'd12479:data <=32'hFFC0FFA3;
14'd12480:data <=32'hFFDCFFA2;14'd12481:data <=32'hFFC9FF8D;14'd12482:data <=32'hFFB3FF90;
14'd12483:data <=32'hFFA0FFCB;14'd12484:data <=32'hFF65FFAE;14'd12485:data <=32'hFF55FFC3;
14'd12486:data <=32'hFF49FFDE;14'd12487:data <=32'hFF44FFFC;14'd12488:data <=32'hFF47001C;
14'd12489:data <=32'hFF54003A;14'd12490:data <=32'hFF680052;14'd12491:data <=32'hFF810061;
14'd12492:data <=32'hFF970067;14'd12493:data <=32'hFFAA0068;14'd12494:data <=32'hFFB70065;
14'd12495:data <=32'hFFBF0062;14'd12496:data <=32'hFFC60064;14'd12497:data <=32'hFFCB0066;
14'd12498:data <=32'hFFD2006C;14'd12499:data <=32'hFFDC0071;14'd12500:data <=32'hFFE90075;
14'd12501:data <=32'hFFF60076;14'd12502:data <=32'h00030076;14'd12503:data <=32'h000F0074;
14'd12504:data <=32'h001D0072;14'd12505:data <=32'h002B006E;14'd12506:data <=32'h003B0067;
14'd12507:data <=32'h004B005C;14'd12508:data <=32'h0059004A;14'd12509:data <=32'h00610033;
14'd12510:data <=32'h00620019;14'd12511:data <=32'h00590001;14'd12512:data <=32'h0047FFED;
14'd12513:data <=32'h002FFFE1;14'd12514:data <=32'h0014FFE0;14'd12515:data <=32'hFFFCFFE9;
14'd12516:data <=32'hFFEAFFFB;14'd12517:data <=32'hFFE00013;14'd12518:data <=32'hFFE1002C;
14'd12519:data <=32'hFFE90043;14'd12520:data <=32'hFFF80058;14'd12521:data <=32'h000D0066;
14'd12522:data <=32'h0025006E;14'd12523:data <=32'h00400071;14'd12524:data <=32'h005C006E;
14'd12525:data <=32'h00780064;14'd12526:data <=32'h00910052;14'd12527:data <=32'h00A70038;
14'd12528:data <=32'h00B6001A;14'd12529:data <=32'h00BBFFF8;14'd12530:data <=32'h00B9FFD6;
14'd12531:data <=32'h00ADFFB8;14'd12532:data <=32'h009CFFA0;14'd12533:data <=32'h0089FF8F;
14'd12534:data <=32'h0076FF83;14'd12535:data <=32'h0069FF7B;14'd12536:data <=32'h005CFF74;
14'd12537:data <=32'h0051FF69;14'd12538:data <=32'h0045FF5E;14'd12539:data <=32'h0035FF4F;
14'd12540:data <=32'h001FFF43;14'd12541:data <=32'h0004FF3A;14'd12542:data <=32'hFFE6FF37;
14'd12543:data <=32'hFFC8FF3B;14'd12544:data <=32'h0015FFE1;14'd12545:data <=32'h0025FFC3;
14'd12546:data <=32'h001AFF9B;14'd12547:data <=32'hFF93FF5E;14'd12548:data <=32'hFF4CFF51;
14'd12549:data <=32'hFF36FF78;14'd12550:data <=32'hFF26FFA4;14'd12551:data <=32'hFF22FFD1;
14'd12552:data <=32'hFF2CFFFD;14'd12553:data <=32'hFF410025;14'd12554:data <=32'hFF5F0042;
14'd12555:data <=32'hFF830052;14'd12556:data <=32'hFFA60054;14'd12557:data <=32'hFFC3004B;
14'd12558:data <=32'hFFD6003A;14'd12559:data <=32'hFFDF0026;14'd12560:data <=32'hFFDD0016;
14'd12561:data <=32'hFFD5000B;14'd12562:data <=32'hFFCA0006;14'd12563:data <=32'hFFBF0009;
14'd12564:data <=32'hFFB5000E;14'd12565:data <=32'hFFAD0018;14'd12566:data <=32'hFFA70024;
14'd12567:data <=32'hFFA50034;14'd12568:data <=32'hFFA70046;14'd12569:data <=32'hFFAF0059;
14'd12570:data <=32'hFFBC006A;14'd12571:data <=32'hFFD00078;14'd12572:data <=32'hFFEA007D;
14'd12573:data <=32'h0003007B;14'd12574:data <=32'h001B0070;14'd12575:data <=32'h002D005E;
14'd12576:data <=32'h00350048;14'd12577:data <=32'h00350034;14'd12578:data <=32'h002F0022;
14'd12579:data <=32'h00220019;14'd12580:data <=32'h00160014;14'd12581:data <=32'h000C0015;
14'd12582:data <=32'h0003001A;14'd12583:data <=32'hFFFF0020;14'd12584:data <=32'hFFFD0026;
14'd12585:data <=32'hFFFB002C;14'd12586:data <=32'hFFFA0033;14'd12587:data <=32'hFFFC003C;
14'd12588:data <=32'hFFFE0046;14'd12589:data <=32'h00030050;14'd12590:data <=32'h000D005A;
14'd12591:data <=32'h001A0063;14'd12592:data <=32'h002B0069;14'd12593:data <=32'h003C006B;
14'd12594:data <=32'h004F006A;14'd12595:data <=32'h00600067;14'd12596:data <=32'h00720062;
14'd12597:data <=32'h0085005B;14'd12598:data <=32'h009B0053;14'd12599:data <=32'h00B50044;
14'd12600:data <=32'h00CF002F;14'd12601:data <=32'h00E70010;14'd12602:data <=32'h00FAFFE5;
14'd12603:data <=32'h0102FFB2;14'd12604:data <=32'h00FAFF7C;14'd12605:data <=32'h00E4FF46;
14'd12606:data <=32'h00BFFF18;14'd12607:data <=32'h0090FEF4;14'd12608:data <=32'h0024FFBC;
14'd12609:data <=32'h0035FFAD;14'd12610:data <=32'h004DFF8B;14'd12611:data <=32'h0051FEFA;
14'd12612:data <=32'hFFEFFECF;14'd12613:data <=32'hFFB6FEE2;14'd12614:data <=32'hFF84FEFF;
14'd12615:data <=32'hFF5CFF26;14'd12616:data <=32'hFF3FFF58;14'd12617:data <=32'hFF34FF8D;
14'd12618:data <=32'hFF37FFBF;14'd12619:data <=32'hFF49FFE8;14'd12620:data <=32'hFF620007;
14'd12621:data <=32'hFF7E0018;14'd12622:data <=32'hFF98001D;14'd12623:data <=32'hFFAC001B;
14'd12624:data <=32'hFFB90015;14'd12625:data <=32'hFFC10010;14'd12626:data <=32'hFFC4000C;
14'd12627:data <=32'hFFC60009;14'd12628:data <=32'hFFC70008;14'd12629:data <=32'hFFC70006;
14'd12630:data <=32'hFFC50004;14'd12631:data <=32'hFFC30004;14'd12632:data <=32'hFFBE0006;
14'd12633:data <=32'hFFB9000C;14'd12634:data <=32'hFFB60014;14'd12635:data <=32'hFFB7001E;
14'd12636:data <=32'hFFBA0027;14'd12637:data <=32'hFFC2002E;14'd12638:data <=32'hFFCA0032;
14'd12639:data <=32'hFFD10032;14'd12640:data <=32'hFFD60031;14'd12641:data <=32'hFFD6002E;
14'd12642:data <=32'hFFD4002E;14'd12643:data <=32'hFFD20034;14'd12644:data <=32'hFFD1003C;
14'd12645:data <=32'hFFD60045;14'd12646:data <=32'hFFDE004E;14'd12647:data <=32'hFFEA0054;
14'd12648:data <=32'hFFF80055;14'd12649:data <=32'h0005004F;14'd12650:data <=32'h000E0046;
14'd12651:data <=32'h0012003B;14'd12652:data <=32'h00100032;14'd12653:data <=32'h000B002B;
14'd12654:data <=32'h00030027;14'd12655:data <=32'hFFF90029;14'd12656:data <=32'hFFF1002F;
14'd12657:data <=32'hFFEB0039;14'd12658:data <=32'hFFE60046;14'd12659:data <=32'hFFE40057;
14'd12660:data <=32'hFFE8006C;14'd12661:data <=32'hFFF20084;14'd12662:data <=32'h0005009D;
14'd12663:data <=32'h002500B3;14'd12664:data <=32'h004E00C1;14'd12665:data <=32'h007F00C3;
14'd12666:data <=32'h00B400B4;14'd12667:data <=32'h00E50095;14'd12668:data <=32'h010D0067;
14'd12669:data <=32'h0127002F;14'd12670:data <=32'h0130FFF1;14'd12671:data <=32'h012BFFB4;
14'd12672:data <=32'h00B7FFDF;14'd12673:data <=32'h00CAFFBF;14'd12674:data <=32'h00DDFFAB;
14'd12675:data <=32'h0100FFA3;14'd12676:data <=32'h00BEFF52;14'd12677:data <=32'h009AFF3A;
14'd12678:data <=32'h0073FF29;14'd12679:data <=32'h004CFF20;14'd12680:data <=32'h0024FF23;
14'd12681:data <=32'h0002FF2E;14'd12682:data <=32'hFFE7FF3E;14'd12683:data <=32'hFFD3FF51;
14'd12684:data <=32'hFFC6FF61;14'd12685:data <=32'hFFBCFF6F;14'd12686:data <=32'hFFB2FF78;
14'd12687:data <=32'hFFA7FF81;14'd12688:data <=32'hFF98FF8C;14'd12689:data <=32'hFF8BFF9C;
14'd12690:data <=32'hFF7FFFB0;14'd12691:data <=32'hFF78FFC9;14'd12692:data <=32'hFF78FFE2;
14'd12693:data <=32'hFF80FFFA;14'd12694:data <=32'hFF8D000E;14'd12695:data <=32'hFF9D001D;
14'd12696:data <=32'hFFAE0025;14'd12697:data <=32'hFFBF0028;14'd12698:data <=32'hFFCF0028;
14'd12699:data <=32'hFFDC0025;14'd12700:data <=32'hFFE9001E;14'd12701:data <=32'hFFF30014;
14'd12702:data <=32'hFFFA0006;14'd12703:data <=32'hFFFAFFF5;14'd12704:data <=32'hFFF4FFE5;
14'd12705:data <=32'hFFE6FFD8;14'd12706:data <=32'hFFD2FFD1;14'd12707:data <=32'hFFBAFFD4;
14'd12708:data <=32'hFFA6FFDE;14'd12709:data <=32'hFF96FFF2;14'd12710:data <=32'hFF8E0008;
14'd12711:data <=32'hFF8F0021;14'd12712:data <=32'hFF980038;14'd12713:data <=32'hFFA60047;
14'd12714:data <=32'hFFB70051;14'd12715:data <=32'hFFC60054;14'd12716:data <=32'hFFD40053;
14'd12717:data <=32'hFFDD0050;14'd12718:data <=32'hFFE3004B;14'd12719:data <=32'hFFE60047;
14'd12720:data <=32'hFFE70044;14'd12721:data <=32'hFFE60043;14'd12722:data <=32'hFFE30044;
14'd12723:data <=32'hFFDF0047;14'd12724:data <=32'hFFD90050;14'd12725:data <=32'hFFD6005D;
14'd12726:data <=32'hFFD60070;14'd12727:data <=32'hFFDE0087;14'd12728:data <=32'hFFF0009D;
14'd12729:data <=32'h000C00B0;14'd12730:data <=32'h002E00BB;14'd12731:data <=32'h005700BA;
14'd12732:data <=32'h007C00AD;14'd12733:data <=32'h009D0095;14'd12734:data <=32'h00B60078;
14'd12735:data <=32'h00C60057;14'd12736:data <=32'h00B800B3;14'd12737:data <=32'h00F3009B;
14'd12738:data <=32'h010E0077;14'd12739:data <=32'h00B1004D;14'd12740:data <=32'h00900011;
14'd12741:data <=32'h00920006;14'd12742:data <=32'h0093FFFB;14'd12743:data <=32'h0095FFED;
14'd12744:data <=32'h0096FFE0;14'd12745:data <=32'h0096FFD2;14'd12746:data <=32'h0096FFC3;
14'd12747:data <=32'h0097FFB1;14'd12748:data <=32'h0095FF9B;14'd12749:data <=32'h0090FF81;
14'd12750:data <=32'h0083FF63;14'd12751:data <=32'h006BFF45;14'd12752:data <=32'h0048FF2D;
14'd12753:data <=32'h001EFF1F;14'd12754:data <=32'hFFEFFF1F;14'd12755:data <=32'hFFC2FF2D;
14'd12756:data <=32'hFF9BFF45;14'd12757:data <=32'hFF7EFF67;14'd12758:data <=32'hFF6DFF8E;
14'd12759:data <=32'hFF67FFB3;14'd12760:data <=32'hFF6BFFD7;14'd12761:data <=32'hFF75FFF7;
14'd12762:data <=32'hFF870011;14'd12763:data <=32'hFF9D0026;14'd12764:data <=32'hFFB70034;
14'd12765:data <=32'hFFD40038;14'd12766:data <=32'hFFEF0034;14'd12767:data <=32'h00080025;
14'd12768:data <=32'h00190011;14'd12769:data <=32'h0022FFF7;14'd12770:data <=32'h001FFFDC;
14'd12771:data <=32'h0013FFC5;14'd12772:data <=32'hFFFFFFB5;14'd12773:data <=32'hFFE9FFAD;
14'd12774:data <=32'hFFD2FFAE;14'd12775:data <=32'hFFC0FFB3;14'd12776:data <=32'hFFB0FFBD;
14'd12777:data <=32'hFFA5FFC7;14'd12778:data <=32'hFF9CFFD1;14'd12779:data <=32'hFF94FFDA;
14'd12780:data <=32'hFF8BFFE4;14'd12781:data <=32'hFF82FFF1;14'd12782:data <=32'hFF790000;
14'd12783:data <=32'hFF730012;14'd12784:data <=32'hFF6F0028;14'd12785:data <=32'hFF71003E;
14'd12786:data <=32'hFF770054;14'd12787:data <=32'hFF810068;14'd12788:data <=32'hFF8C007B;
14'd12789:data <=32'hFF9B008D;14'd12790:data <=32'hFFAB009E;14'd12791:data <=32'hFFC000AD;
14'd12792:data <=32'hFFDA00BA;14'd12793:data <=32'hFFF800C3;14'd12794:data <=32'h001A00C3;
14'd12795:data <=32'h003C00B9;14'd12796:data <=32'h005B00A7;14'd12797:data <=32'h0072008D;
14'd12798:data <=32'h007D006F;14'd12799:data <=32'h007F0052;14'd12800:data <=32'hFFFA00E8;
14'd12801:data <=32'h00310101;14'd12802:data <=32'h006C00F3;14'd12803:data <=32'h006E0052;
14'd12804:data <=32'h00410020;14'd12805:data <=32'h00390027;14'd12806:data <=32'h00370030;
14'd12807:data <=32'h003B003A;14'd12808:data <=32'h00430043;14'd12809:data <=32'h0051004B;
14'd12810:data <=32'h0064004E;14'd12811:data <=32'h007C004B;14'd12812:data <=32'h00970041;
14'd12813:data <=32'h00B1002A;14'd12814:data <=32'h00C50009;14'd12815:data <=32'h00D0FFE0;
14'd12816:data <=32'h00CCFFB4;14'd12817:data <=32'h00BAFF88;14'd12818:data <=32'h009CFF65;
14'd12819:data <=32'h0075FF4C;14'd12820:data <=32'h004CFF41;14'd12821:data <=32'h0024FF40;
14'd12822:data <=32'h0000FF48;14'd12823:data <=32'hFFE2FF58;14'd12824:data <=32'hFFC9FF6B;
14'd12825:data <=32'hFFB7FF82;14'd12826:data <=32'hFFAAFF99;14'd12827:data <=32'hFFA2FFB3;
14'd12828:data <=32'hFFA2FFCE;14'd12829:data <=32'hFFA7FFE6;14'd12830:data <=32'hFFB5FFFB;
14'd12831:data <=32'hFFC6000A;14'd12832:data <=32'hFFDB0011;14'd12833:data <=32'hFFEE0012;
14'd12834:data <=32'hFFFF000B;14'd12835:data <=32'h000B0001;14'd12836:data <=32'h0013FFF6;
14'd12837:data <=32'h0017FFEB;14'd12838:data <=32'h001AFFDF;14'd12839:data <=32'h001CFFD5;
14'd12840:data <=32'h001DFFC8;14'd12841:data <=32'h001CFFB9;14'd12842:data <=32'h0018FFA6;
14'd12843:data <=32'h000CFF91;14'd12844:data <=32'hFFF8FF7C;14'd12845:data <=32'hFFDBFF6C;
14'd12846:data <=32'hFFB8FF65;14'd12847:data <=32'hFF91FF67;14'd12848:data <=32'hFF6AFF75;
14'd12849:data <=32'hFF47FF8E;14'd12850:data <=32'hFF29FFAF;14'd12851:data <=32'hFF15FFD7;
14'd12852:data <=32'hFF0A0003;14'd12853:data <=32'hFF080031;14'd12854:data <=32'hFF0F0060;
14'd12855:data <=32'hFF21008E;14'd12856:data <=32'hFF3E00B7;14'd12857:data <=32'hFF6500DA;
14'd12858:data <=32'hFF9500F3;14'd12859:data <=32'hFFCA00FD;14'd12860:data <=32'hFFFF00F7;
14'd12861:data <=32'h002E00E3;14'd12862:data <=32'h005200C3;14'd12863:data <=32'h0068009E;
14'd12864:data <=32'hFFC10088;14'd12865:data <=32'hFFCF00A4;14'd12866:data <=32'hFFF700C1;
14'd12867:data <=32'h005D00A5;14'd12868:data <=32'h003E0065;14'd12869:data <=32'h003D005D;
14'd12870:data <=32'h003C0058;14'd12871:data <=32'h003E0056;14'd12872:data <=32'h00400055;
14'd12873:data <=32'h00430054;14'd12874:data <=32'h004A0055;14'd12875:data <=32'h00540056;
14'd12876:data <=32'h00610054;14'd12877:data <=32'h0073004E;14'd12878:data <=32'h00840041;
14'd12879:data <=32'h0093002C;14'd12880:data <=32'h009B0012;14'd12881:data <=32'h009AFFF7;
14'd12882:data <=32'h0091FFDD;14'd12883:data <=32'h0081FFC9;14'd12884:data <=32'h006FFFBC;
14'd12885:data <=32'h005DFFB5;14'd12886:data <=32'h0050FFB4;14'd12887:data <=32'h0045FFB4;
14'd12888:data <=32'h003CFFB3;14'd12889:data <=32'h0035FFB1;14'd12890:data <=32'h002DFFAE;
14'd12891:data <=32'h0024FFAC;14'd12892:data <=32'h0018FFAB;14'd12893:data <=32'h000CFFAF;
14'd12894:data <=32'h0004FFB2;14'd12895:data <=32'hFFFBFFB9;14'd12896:data <=32'hFFF7FFC0;
14'd12897:data <=32'hFFF1FFC6;14'd12898:data <=32'hFFEEFFCE;14'd12899:data <=32'hFFECFFD5;
14'd12900:data <=32'hFFEBFFDF;14'd12901:data <=32'hFFECFFE9;14'd12902:data <=32'hFFF2FFF5;
14'd12903:data <=32'hFFFEFFFF;14'd12904:data <=32'h000F0005;14'd12905:data <=32'h00250003;
14'd12906:data <=32'h003BFFF6;14'd12907:data <=32'h004DFFE0;14'd12908:data <=32'h0059FFC2;
14'd12909:data <=32'h0058FF9F;14'd12910:data <=32'h004AFF7A;14'd12911:data <=32'h0030FF5A;
14'd12912:data <=32'h000DFF42;14'd12913:data <=32'hFFE4FF34;14'd12914:data <=32'hFFB8FF32;
14'd12915:data <=32'hFF8CFF3A;14'd12916:data <=32'hFF63FF4B;14'd12917:data <=32'hFF3DFF66;
14'd12918:data <=32'hFF1EFF8A;14'd12919:data <=32'hFF06FFB4;14'd12920:data <=32'hFEF8FFE4;
14'd12921:data <=32'hFEF60017;14'd12922:data <=32'hFF020049;14'd12923:data <=32'hFF1A0075;
14'd12924:data <=32'hFF3C0097;14'd12925:data <=32'hFF6200AD;14'd12926:data <=32'hFF8800B7;
14'd12927:data <=32'hFFA900B7;14'd12928:data <=32'hFFBB0094;14'd12929:data <=32'hFFC6009C;
14'd12930:data <=32'hFFC800AE;14'd12931:data <=32'hFF9C00D4;14'd12932:data <=32'hFF9400B2;
14'd12933:data <=32'hFFAB00C4;14'd12934:data <=32'hFFCA00D1;14'd12935:data <=32'hFFEC00D9;
14'd12936:data <=32'h000E00D8;14'd12937:data <=32'h003000D0;14'd12938:data <=32'h004D00C1;
14'd12939:data <=32'h006700AF;14'd12940:data <=32'h007E0099;14'd12941:data <=32'h00920080;
14'd12942:data <=32'h00A10062;14'd12943:data <=32'h00A80041;14'd12944:data <=32'h00A7001C;
14'd12945:data <=32'h009BFFFB;14'd12946:data <=32'h0087FFE0;14'd12947:data <=32'h006BFFCE;
14'd12948:data <=32'h004EFFC8;14'd12949:data <=32'h0033FFCC;14'd12950:data <=32'h0020FFDB;
14'd12951:data <=32'h0017FFEC;14'd12952:data <=32'h0016FFFD;14'd12953:data <=32'h001C0008;
14'd12954:data <=32'h0026000F;14'd12955:data <=32'h0031000F;14'd12956:data <=32'h003B000D;
14'd12957:data <=32'h00420007;14'd12958:data <=32'h0049FFFF;14'd12959:data <=32'h004CFFF5;
14'd12960:data <=32'h004DFFEA;14'd12961:data <=32'h004CFFDE;14'd12962:data <=32'h0047FFD2;
14'd12963:data <=32'h003DFFC8;14'd12964:data <=32'h0031FFC2;14'd12965:data <=32'h0023FFC1;
14'd12966:data <=32'h0016FFC7;14'd12967:data <=32'h000EFFD1;14'd12968:data <=32'h000CFFDE;
14'd12969:data <=32'h0012FFE9;14'd12970:data <=32'h001FFFF1;14'd12971:data <=32'h002FFFF0;
14'd12972:data <=32'h003EFFE8;14'd12973:data <=32'h004BFFD7;14'd12974:data <=32'h0050FFC2;
14'd12975:data <=32'h004EFFAC;14'd12976:data <=32'h0046FF96;14'd12977:data <=32'h0037FF84;
14'd12978:data <=32'h0026FF76;14'd12979:data <=32'h0012FF6C;14'd12980:data <=32'hFFFDFF65;
14'd12981:data <=32'hFFE8FF5F;14'd12982:data <=32'hFFD0FF5F;14'd12983:data <=32'hFFB9FF61;
14'd12984:data <=32'hFF9FFF69;14'd12985:data <=32'hFF89FF74;14'd12986:data <=32'hFF75FF85;
14'd12987:data <=32'hFF66FF99;14'd12988:data <=32'hFF5BFFAD;14'd12989:data <=32'hFF52FFBF;
14'd12990:data <=32'hFF4CFFD0;14'd12991:data <=32'hFF43FFE0;14'd12992:data <=32'hFF42005A;
14'd12993:data <=32'hFF4C006F;14'd12994:data <=32'hFF55006E;14'd12995:data <=32'hFF180006;
14'd12996:data <=32'hFEECFFFF;14'd12997:data <=32'hFEE60036;14'd12998:data <=32'hFEEF0070;
14'd12999:data <=32'hFF0700A7;14'd13000:data <=32'hFF2D00D4;14'd13001:data <=32'hFF5B00F5;
14'd13002:data <=32'hFF8F010C;14'd13003:data <=32'hFFC50116;14'd13004:data <=32'hFFFB0116;
14'd13005:data <=32'h00300109;14'd13006:data <=32'h006000F0;14'd13007:data <=32'h008800CD;
14'd13008:data <=32'h00A6009F;14'd13009:data <=32'h00B4006D;14'd13010:data <=32'h00B3003A;
14'd13011:data <=32'h00A30010;14'd13012:data <=32'h0088FFEE;14'd13013:data <=32'h0069FFDA;
14'd13014:data <=32'h0048FFD3;14'd13015:data <=32'h002DFFD8;14'd13016:data <=32'h0019FFE2;
14'd13017:data <=32'h000CFFEF;14'd13018:data <=32'h0006FFFD;14'd13019:data <=32'h0004000A;
14'd13020:data <=32'h00040014;14'd13021:data <=32'h0008001F;14'd13022:data <=32'h000D0028;
14'd13023:data <=32'h0016002F;14'd13024:data <=32'h00200035;14'd13025:data <=32'h002D0035;
14'd13026:data <=32'h003A0034;14'd13027:data <=32'h0046002D;14'd13028:data <=32'h004F0024;
14'd13029:data <=32'h0055001A;14'd13030:data <=32'h00570011;14'd13031:data <=32'h005A000A;
14'd13032:data <=32'h005D0003;14'd13033:data <=32'h0060FFFD;14'd13034:data <=32'h0066FFF5;
14'd13035:data <=32'h006CFFE9;14'd13036:data <=32'h0070FFDA;14'd13037:data <=32'h0070FFC6;
14'd13038:data <=32'h006AFFB2;14'd13039:data <=32'h005CFF9F;14'd13040:data <=32'h004AFF92;
14'd13041:data <=32'h0036FF8C;14'd13042:data <=32'h0022FF8D;14'd13043:data <=32'h0012FF91;
14'd13044:data <=32'h0008FF9B;14'd13045:data <=32'h0002FFA3;14'd13046:data <=32'h0001FFAA;
14'd13047:data <=32'h0003FFAD;14'd13048:data <=32'h0005FFAC;14'd13049:data <=32'h0006FFA8;
14'd13050:data <=32'h0008FFA2;14'd13051:data <=32'h0007FF99;14'd13052:data <=32'h0004FF8C;
14'd13053:data <=32'hFFFEFF7C;14'd13054:data <=32'hFFF1FF69;14'd13055:data <=32'hFFDBFF55;
14'd13056:data <=32'hFF6CFF92;14'd13057:data <=32'hFF55FF99;14'd13058:data <=32'hFF56FFA4;
14'd13059:data <=32'hFF99FF64;14'd13060:data <=32'hFF51FF3F;14'd13061:data <=32'hFF24FF5F;
14'd13062:data <=32'hFF03FF8D;14'd13063:data <=32'hFEEFFFC2;14'd13064:data <=32'hFEE9FFF8;
14'd13065:data <=32'hFEF0002B;14'd13066:data <=32'hFEFF005A;14'd13067:data <=32'hFF190085;
14'd13068:data <=32'hFF3800A8;14'd13069:data <=32'hFF6000C5;14'd13070:data <=32'hFF8C00D7;
14'd13071:data <=32'hFFBA00DF;14'd13072:data <=32'hFFE800DA;14'd13073:data <=32'h001100CA;
14'd13074:data <=32'h003000B0;14'd13075:data <=32'h00450093;14'd13076:data <=32'h004F0075;
14'd13077:data <=32'h0051005C;14'd13078:data <=32'h004E0048;14'd13079:data <=32'h00490039;
14'd13080:data <=32'h0046002D;14'd13081:data <=32'h00430023;14'd13082:data <=32'h003E0018;
14'd13083:data <=32'h0039000D;14'd13084:data <=32'h002F0003;14'd13085:data <=32'h0023FFFB;
14'd13086:data <=32'h0014FFF8;14'd13087:data <=32'h0004FFFC;14'd13088:data <=32'hFFF60004;
14'd13089:data <=32'hFFED0012;14'd13090:data <=32'hFFE80021;14'd13091:data <=32'hFFE90031;
14'd13092:data <=32'hFFEE0042;14'd13093:data <=32'hFFF80051;14'd13094:data <=32'h0005005E;
14'd13095:data <=32'h00160069;14'd13096:data <=32'h002B0071;14'd13097:data <=32'h00440076;
14'd13098:data <=32'h00620072;14'd13099:data <=32'h007F0066;14'd13100:data <=32'h009B004F;
14'd13101:data <=32'h00AF0030;14'd13102:data <=32'h00BB000B;14'd13103:data <=32'h00BBFFE5;
14'd13104:data <=32'h00AEFFC0;14'd13105:data <=32'h0098FFA3;14'd13106:data <=32'h007CFF91;
14'd13107:data <=32'h005FFF88;14'd13108:data <=32'h0045FF88;14'd13109:data <=32'h0030FF8E;
14'd13110:data <=32'h0023FF97;14'd13111:data <=32'h001AFFA1;14'd13112:data <=32'h0016FFAA;
14'd13113:data <=32'h0016FFB2;14'd13114:data <=32'h0019FFB7;14'd13115:data <=32'h001FFFB9;
14'd13116:data <=32'h0027FFB5;14'd13117:data <=32'h0031FFAB;14'd13118:data <=32'h0036FF9A;
14'd13119:data <=32'h0035FF82;14'd13120:data <=32'h0037FF89;14'd13121:data <=32'h002DFF63;
14'd13122:data <=32'h0017FF54;14'd13123:data <=32'hFFF7FF7D;14'd13124:data <=32'hFFC1FF45;
14'd13125:data <=32'hFF9FFF51;14'd13126:data <=32'hFF84FF66;14'd13127:data <=32'hFF6FFF81;
14'd13128:data <=32'hFF63FF9C;14'd13129:data <=32'hFF5DFFB6;14'd13130:data <=32'hFF5DFFCC;
14'd13131:data <=32'hFF5DFFE1;14'd13132:data <=32'hFF5FFFF3;14'd13133:data <=32'hFF620007;
14'd13134:data <=32'hFF68001A;14'd13135:data <=32'hFF71002A;14'd13136:data <=32'hFF7D0038;
14'd13137:data <=32'hFF8A0043;14'd13138:data <=32'hFF96004A;14'd13139:data <=32'hFF9F0050;
14'd13140:data <=32'hFFA60055;14'd13141:data <=32'hFFAD005D;14'd13142:data <=32'hFFB40068;
14'd13143:data <=32'hFFC20074;14'd13144:data <=32'hFFD4007E;14'd13145:data <=32'hFFEC0084;
14'd13146:data <=32'h00060082;14'd13147:data <=32'h001F0077;14'd13148:data <=32'h00340063;
14'd13149:data <=32'h00400049;14'd13150:data <=32'h00430030;14'd13151:data <=32'h003D0018;
14'd13152:data <=32'h002F0004;14'd13153:data <=32'h001DFFF8;14'd13154:data <=32'h0009FFF2;
14'd13155:data <=32'hFFF5FFF3;14'd13156:data <=32'hFFE2FFFB;14'd13157:data <=32'hFFD10007;
14'd13158:data <=32'hFFC4001A;14'd13159:data <=32'hFFBD0031;14'd13160:data <=32'hFFBD004D;
14'd13161:data <=32'hFFC60069;14'd13162:data <=32'hFFD90083;14'd13163:data <=32'hFFF50097;
14'd13164:data <=32'h001700A3;14'd13165:data <=32'h003C00A4;14'd13166:data <=32'h005F0099;
14'd13167:data <=32'h007C0084;14'd13168:data <=32'h0092006B;14'd13169:data <=32'h009E004F;
14'd13170:data <=32'h00A20035;14'd13171:data <=32'h00A3001F;14'd13172:data <=32'h00A1000C;
14'd13173:data <=32'h009EFFFC;14'd13174:data <=32'h009DFFED;14'd13175:data <=32'h009BFFDD;
14'd13176:data <=32'h0099FFCC;14'd13177:data <=32'h0093FFBB;14'd13178:data <=32'h008CFFAA;
14'd13179:data <=32'h0082FF9A;14'd13180:data <=32'h0078FF8C;14'd13181:data <=32'h006DFF7F;
14'd13182:data <=32'h0061FF72;14'd13183:data <=32'h0054FF62;14'd13184:data <=32'h005A000B;
14'd13185:data <=32'h0080FFE9;14'd13186:data <=32'h0086FFB5;14'd13187:data <=32'h0018FF4D;
14'd13188:data <=32'hFFD9FF1D;14'd13189:data <=32'hFFB1FF34;14'd13190:data <=32'hFF94FF53;
14'd13191:data <=32'hFF81FF78;14'd13192:data <=32'hFF7CFF9E;14'd13193:data <=32'hFF83FFBD;
14'd13194:data <=32'hFF90FFD5;14'd13195:data <=32'hFFA1FFE3;14'd13196:data <=32'hFFB0FFE9;
14'd13197:data <=32'hFFBCFFE9;14'd13198:data <=32'hFFC4FFE7;14'd13199:data <=32'hFFC9FFE2;
14'd13200:data <=32'hFFCBFFDC;14'd13201:data <=32'hFFCAFFD5;14'd13202:data <=32'hFFC2FFCE;
14'd13203:data <=32'hFFB6FFC9;14'd13204:data <=32'hFFA4FFC9;14'd13205:data <=32'hFF91FFD0;
14'd13206:data <=32'hFF7EFFE1;14'd13207:data <=32'hFF71FFFA;14'd13208:data <=32'hFF6D0017;
14'd13209:data <=32'hFF740038;14'd13210:data <=32'hFF860053;14'd13211:data <=32'hFF9D0067;
14'd13212:data <=32'hFFBA0070;14'd13213:data <=32'hFFD6006F;14'd13214:data <=32'hFFEE0068;
14'd13215:data <=32'h0000005A;14'd13216:data <=32'h000B004B;14'd13217:data <=32'h0012003B;
14'd13218:data <=32'h0013002C;14'd13219:data <=32'h0010001E;14'd13220:data <=32'h000A0012;
14'd13221:data <=32'h00010009;14'd13222:data <=32'hFFF40002;14'd13223:data <=32'hFFE60001;
14'd13224:data <=32'hFFD60006;14'd13225:data <=32'hFFC80010;14'd13226:data <=32'hFFBE0020;
14'd13227:data <=32'hFFB90033;14'd13228:data <=32'hFFBB0047;14'd13229:data <=32'hFFC20058;
14'd13230:data <=32'hFFCD0067;14'd13231:data <=32'hFFDA0071;14'd13232:data <=32'hFFE6007B;
14'd13233:data <=32'hFFF10083;14'd13234:data <=32'hFFFD008D;14'd13235:data <=32'h000C0099;
14'd13236:data <=32'h002000A6;14'd13237:data <=32'h003A00B1;14'd13238:data <=32'h005C00B6;
14'd13239:data <=32'h008200B1;14'd13240:data <=32'h00A900A3;14'd13241:data <=32'h00CE0089;
14'd13242:data <=32'h00ED0066;14'd13243:data <=32'h0103003B;14'd13244:data <=32'h010F000D;
14'd13245:data <=32'h0113FFDC;14'd13246:data <=32'h010CFFAC;14'd13247:data <=32'h00FCFF7C;
14'd13248:data <=32'h00480010;14'd13249:data <=32'h006E000A;14'd13250:data <=32'h009CFFEA;
14'd13251:data <=32'h00CEFF4F;14'd13252:data <=32'h0085FEFB;14'd13253:data <=32'h0049FEF6;
14'd13254:data <=32'h000EFF00;14'd13255:data <=32'hFFDFFF18;14'd13256:data <=32'hFFBCFF3B;
14'd13257:data <=32'hFFA8FF61;14'd13258:data <=32'hFFA1FF83;14'd13259:data <=32'hFFA3FFA1;
14'd13260:data <=32'hFFA9FFB8;14'd13261:data <=32'hFFB2FFC8;14'd13262:data <=32'hFFBDFFD3;
14'd13263:data <=32'hFFC9FFDA;14'd13264:data <=32'hFFD3FFDD;14'd13265:data <=32'hFFDCFFDC;
14'd13266:data <=32'hFFE4FFD5;14'd13267:data <=32'hFFE6FFCC;14'd13268:data <=32'hFFE1FFC2;
14'd13269:data <=32'hFFD6FFBA;14'd13270:data <=32'hFFC7FFB7;14'd13271:data <=32'hFFB5FFBC;
14'd13272:data <=32'hFFA8FFC7;14'd13273:data <=32'hFF9EFFD7;14'd13274:data <=32'hFF9CFFE9;
14'd13275:data <=32'hFF9FFFF9;14'd13276:data <=32'hFFA60005;14'd13277:data <=32'hFFAF000C;
14'd13278:data <=32'hFFB6000F;14'd13279:data <=32'hFFBA0011;14'd13280:data <=32'hFFBD0012;
14'd13281:data <=32'hFFBC0016;14'd13282:data <=32'hFFBE001B;14'd13283:data <=32'hFFC10021;
14'd13284:data <=32'hFFC70027;14'd13285:data <=32'hFFCD002A;14'd13286:data <=32'hFFD5002B;
14'd13287:data <=32'hFFDB0029;14'd13288:data <=32'hFFE00027;14'd13289:data <=32'hFFE20022;
14'd13290:data <=32'hFFE3001F;14'd13291:data <=32'hFFE2001C;14'd13292:data <=32'hFFE00018;
14'd13293:data <=32'hFFDC0016;14'd13294:data <=32'hFFD70012;14'd13295:data <=32'hFFCE000F;
14'd13296:data <=32'hFFC1000F;14'd13297:data <=32'hFFAF0015;14'd13298:data <=32'hFF9C0024;
14'd13299:data <=32'hFF8B003C;14'd13300:data <=32'hFF83005F;14'd13301:data <=32'hFF840089;
14'd13302:data <=32'hFF9500B2;14'd13303:data <=32'hFFB300D9;14'd13304:data <=32'hFFDF00F7;
14'd13305:data <=32'h00130109;14'd13306:data <=32'h004B010D;14'd13307:data <=32'h00830103;
14'd13308:data <=32'h00B700EB;14'd13309:data <=32'h00E500C9;14'd13310:data <=32'h010C009C;
14'd13311:data <=32'h01290068;14'd13312:data <=32'h00990056;14'd13313:data <=32'h00C00048;
14'd13314:data <=32'h00E50040;14'd13315:data <=32'h01210038;14'd13316:data <=32'h0104FFCC;
14'd13317:data <=32'h00EAFFA4;14'd13318:data <=32'h00CAFF87;14'd13319:data <=32'h00A7FF74;
14'd13320:data <=32'h0088FF6B;14'd13321:data <=32'h006EFF69;14'd13322:data <=32'h0058FF68;
14'd13323:data <=32'h0047FF68;14'd13324:data <=32'h0036FF66;14'd13325:data <=32'h0023FF65;
14'd13326:data <=32'h0010FF65;14'd13327:data <=32'hFFFDFF6A;14'd13328:data <=32'hFFE9FF74;
14'd13329:data <=32'hFFDAFF80;14'd13330:data <=32'hFFCFFF8C;14'd13331:data <=32'hFFC6FF99;
14'd13332:data <=32'hFFBFFFA5;14'd13333:data <=32'hFFBAFFB2;14'd13334:data <=32'hFFB6FFBE;
14'd13335:data <=32'hFFB2FFCD;14'd13336:data <=32'hFFB3FFDD;14'd13337:data <=32'hFFB8FFED;
14'd13338:data <=32'hFFC5FFFB;14'd13339:data <=32'hFFD40002;14'd13340:data <=32'hFFE50002;
14'd13341:data <=32'hFFF4FFF9;14'd13342:data <=32'hFFFDFFEB;14'd13343:data <=32'hFFFEFFDB;
14'd13344:data <=32'hFFF8FFCB;14'd13345:data <=32'hFFEAFFBF;14'd13346:data <=32'hFFD8FFBA;
14'd13347:data <=32'hFFC7FFBD;14'd13348:data <=32'hFFB7FFC5;14'd13349:data <=32'hFFABFFD1;
14'd13350:data <=32'hFFA4FFDF;14'd13351:data <=32'hFFA1FFED;14'd13352:data <=32'hFFA2FFFB;
14'd13353:data <=32'hFFA50007;14'd13354:data <=32'hFFAA0012;14'd13355:data <=32'hFFB20019;
14'd13356:data <=32'hFFBB0020;14'd13357:data <=32'hFFC50020;14'd13358:data <=32'hFFCD001D;
14'd13359:data <=32'hFFD30015;14'd13360:data <=32'hFFD1000A;14'd13361:data <=32'hFFC80000;
14'd13362:data <=32'hFFB8FFFB;14'd13363:data <=32'hFFA1FFFE;14'd13364:data <=32'hFF8B000B;
14'd13365:data <=32'hFF790023;14'd13366:data <=32'hFF6E0043;14'd13367:data <=32'hFF6F0067;
14'd13368:data <=32'hFF7B008C;14'd13369:data <=32'hFF9100AC;14'd13370:data <=32'hFFAF00C5;
14'd13371:data <=32'hFFD100D6;14'd13372:data <=32'hFFF500E1;14'd13373:data <=32'h001A00E4;
14'd13374:data <=32'h004000E1;14'd13375:data <=32'h006500D6;14'd13376:data <=32'h00410106;
14'd13377:data <=32'h0082010D;14'd13378:data <=32'h00AE00FE;14'd13379:data <=32'h007300C5;
14'd13380:data <=32'h00740079;14'd13381:data <=32'h007D006C;14'd13382:data <=32'h00830061;
14'd13383:data <=32'h008B0058;14'd13384:data <=32'h00960050;14'd13385:data <=32'h00A50046;
14'd13386:data <=32'h00B70036;14'd13387:data <=32'h00CA001E;14'd13388:data <=32'h00D6FFFD;
14'd13389:data <=32'h00DBFFD6;14'd13390:data <=32'h00D3FFAD;14'd13391:data <=32'h00C0FF86;
14'd13392:data <=32'h00A4FF65;14'd13393:data <=32'h0081FF4F;14'd13394:data <=32'h005BFF41;
14'd13395:data <=32'h0035FF3B;14'd13396:data <=32'h0010FF3D;14'd13397:data <=32'hFFECFF48;
14'd13398:data <=32'hFFCAFF5A;14'd13399:data <=32'hFFAFFF74;14'd13400:data <=32'hFF9CFF93;
14'd13401:data <=32'hFF93FFB8;14'd13402:data <=32'hFF96FFDC;14'd13403:data <=32'hFFA5FFFD;
14'd13404:data <=32'hFFBE0015;14'd13405:data <=32'hFFDB0020;14'd13406:data <=32'hFFF9001F;
14'd13407:data <=32'h00120014;14'd13408:data <=32'h00230002;14'd13409:data <=32'h002CFFEC;
14'd13410:data <=32'h002CFFD8;14'd13411:data <=32'h0026FFC5;14'd13412:data <=32'h001BFFB6;
14'd13413:data <=32'h000FFFAC;14'd13414:data <=32'h0001FFA5;14'd13415:data <=32'hFFF4FF9F;
14'd13416:data <=32'hFFE5FF9C;14'd13417:data <=32'hFFD5FF9C;14'd13418:data <=32'hFFC5FF9E;
14'd13419:data <=32'hFFB6FFA4;14'd13420:data <=32'hFFA9FFAE;14'd13421:data <=32'hFF9DFFB9;
14'd13422:data <=32'hFF96FFC3;14'd13423:data <=32'hFF90FFCF;14'd13424:data <=32'hFF8BFFD7;
14'd13425:data <=32'hFF84FFE0;14'd13426:data <=32'hFF7CFFE9;14'd13427:data <=32'hFF71FFF5;
14'd13428:data <=32'hFF670007;14'd13429:data <=32'hFF5F001F;14'd13430:data <=32'hFF5E003A;
14'd13431:data <=32'hFF660057;14'd13432:data <=32'hFF760072;14'd13433:data <=32'hFF8C0087;
14'd13434:data <=32'hFFA70093;14'd13435:data <=32'hFFC10098;14'd13436:data <=32'hFFD70096;
14'd13437:data <=32'hFFEA0090;14'd13438:data <=32'hFFF8008A;14'd13439:data <=32'h00020084;
14'd13440:data <=32'hFF6B00DC;14'd13441:data <=32'hFF960112;14'd13442:data <=32'hFFD40120;
14'd13443:data <=32'h0009008B;14'd13444:data <=32'hFFFA004F;14'd13445:data <=32'hFFF20054;
14'd13446:data <=32'hFFEC0062;14'd13447:data <=32'hFFEC0074;14'd13448:data <=32'hFFF5008B;
14'd13449:data <=32'h000900A3;14'd13450:data <=32'h002900B4;14'd13451:data <=32'h005200BA;
14'd13452:data <=32'h007E00B2;14'd13453:data <=32'h00A7009C;14'd13454:data <=32'h00C9007A;
14'd13455:data <=32'h00DE004F;14'd13456:data <=32'h00E90021;14'd13457:data <=32'h00E7FFF5;
14'd13458:data <=32'h00DBFFCB;14'd13459:data <=32'h00C8FFA6;14'd13460:data <=32'h00AEFF86;
14'd13461:data <=32'h008EFF6E;14'd13462:data <=32'h0069FF5D;14'd13463:data <=32'h0042FF57;
14'd13464:data <=32'h001AFF5B;14'd13465:data <=32'hFFF6FF69;14'd13466:data <=32'hFFDAFF81;
14'd13467:data <=32'hFFC9FF9E;14'd13468:data <=32'hFFC3FFBC;14'd13469:data <=32'hFFC7FFD8;
14'd13470:data <=32'hFFD2FFED;14'd13471:data <=32'hFFE0FFFB;14'd13472:data <=32'hFFEE0003;
14'd13473:data <=32'hFFFC0005;14'd13474:data <=32'h00080006;14'd13475:data <=32'h00130006;
14'd13476:data <=32'h001E0004;14'd13477:data <=32'h002BFFFF;14'd13478:data <=32'h0037FFF7;
14'd13479:data <=32'h0044FFEB;14'd13480:data <=32'h004FFFD9;14'd13481:data <=32'h0053FFC2;
14'd13482:data <=32'h0052FFA9;14'd13483:data <=32'h0049FF8F;14'd13484:data <=32'h0039FF77;
14'd13485:data <=32'h0023FF63;14'd13486:data <=32'h0008FF53;14'd13487:data <=32'hFFEBFF49;
14'd13488:data <=32'hFFCAFF45;14'd13489:data <=32'hFFA6FF46;14'd13490:data <=32'hFF81FF4E;
14'd13491:data <=32'hFF5BFF60;14'd13492:data <=32'hFF38FF7D;14'd13493:data <=32'hFF1AFFA3;
14'd13494:data <=32'hFF08FFD2;14'd13495:data <=32'hFF040005;14'd13496:data <=32'hFF0E0038;
14'd13497:data <=32'hFF260064;14'd13498:data <=32'hFF490086;14'd13499:data <=32'hFF70009B;
14'd13500:data <=32'hFF9700A2;14'd13501:data <=32'hFFBA009E;14'd13502:data <=32'hFFD70094;
14'd13503:data <=32'hFFEB0086;14'd13504:data <=32'hFF5C003F;14'd13505:data <=32'hFF580069;
14'd13506:data <=32'hFF720098;14'd13507:data <=32'hFFEA009B;14'd13508:data <=32'hFFE60055;
14'd13509:data <=32'hFFE1004F;14'd13510:data <=32'hFFD9004F;14'd13511:data <=32'hFFD20055;
14'd13512:data <=32'hFFCD0063;14'd13513:data <=32'hFFD00077;14'd13514:data <=32'hFFDC008D;
14'd13515:data <=32'hFFF3009F;14'd13516:data <=32'h000F00A8;14'd13517:data <=32'h002F00A7;
14'd13518:data <=32'h004D009C;14'd13519:data <=32'h0066008C;14'd13520:data <=32'h00790076;
14'd13521:data <=32'h0084005E;14'd13522:data <=32'h008B0049;14'd13523:data <=32'h008F0033;
14'd13524:data <=32'h0090001E;14'd13525:data <=32'h008E000A;14'd13526:data <=32'h0088FFF6;
14'd13527:data <=32'h007EFFE3;14'd13528:data <=32'h0071FFD4;14'd13529:data <=32'h0061FFCA;
14'd13530:data <=32'h0051FFC3;14'd13531:data <=32'h0043FFC2;14'd13532:data <=32'h0036FFC4;
14'd13533:data <=32'h002EFFC7;14'd13534:data <=32'h0027FFC8;14'd13535:data <=32'h0022FFC8;
14'd13536:data <=32'h0019FFC8;14'd13537:data <=32'h000FFFCA;14'd13538:data <=32'h0003FFCF;
14'd13539:data <=32'hFFF9FFD9;14'd13540:data <=32'hFFF3FFEA;14'd13541:data <=32'hFFF3FFFC;
14'd13542:data <=32'hFFFC000F;14'd13543:data <=32'h000D001F;14'd13544:data <=32'h00250027;
14'd13545:data <=32'h00410026;14'd13546:data <=32'h005B001B;14'd13547:data <=32'h00720007;
14'd13548:data <=32'h0084FFEC;14'd13549:data <=32'h008FFFCC;14'd13550:data <=32'h0090FFA9;
14'd13551:data <=32'h0089FF84;14'd13552:data <=32'h0079FF60;14'd13553:data <=32'h0060FF3D;
14'd13554:data <=32'h003CFF20;14'd13555:data <=32'h000FFF0B;14'd13556:data <=32'hFFDCFF02;
14'd13557:data <=32'hFFA6FF08;14'd13558:data <=32'hFF73FF1C;14'd13559:data <=32'hFF48FF3F;
14'd13560:data <=32'hFF28FF6A;14'd13561:data <=32'hFF18FF9A;14'd13562:data <=32'hFF15FFC8;
14'd13563:data <=32'hFF1DFFF1;14'd13564:data <=32'hFF2B0012;14'd13565:data <=32'hFF3D002C;
14'd13566:data <=32'hFF50003E;14'd13567:data <=32'hFF62004D;14'd13568:data <=32'hFF82002F;
14'd13569:data <=32'hFF80003C;14'd13570:data <=32'hFF760052;14'd13571:data <=32'hFF4B0076;
14'd13572:data <=32'hFF520050;14'd13573:data <=32'hFF5E0064;14'd13574:data <=32'hFF6B0075;
14'd13575:data <=32'hFF7B0087;14'd13576:data <=32'hFF8C0098;14'd13577:data <=32'hFFA100AA;
14'd13578:data <=32'hFFBD00B7;14'd13579:data <=32'hFFDD00C0;14'd13580:data <=32'h000100C0;
14'd13581:data <=32'h002500B5;14'd13582:data <=32'h0041009F;14'd13583:data <=32'h00550083;
14'd13584:data <=32'h005F0065;14'd13585:data <=32'h005E004A;14'd13586:data <=32'h00560034;
14'd13587:data <=32'h004B0025;14'd13588:data <=32'h003E001D;14'd13589:data <=32'h0034001B;
14'd13590:data <=32'h002D001B;14'd13591:data <=32'h0027001D;14'd13592:data <=32'h00240021;
14'd13593:data <=32'h00230026;14'd13594:data <=32'h0025002A;14'd13595:data <=32'h002B0030;
14'd13596:data <=32'h00330032;14'd13597:data <=32'h003F0032;14'd13598:data <=32'h004C002B;
14'd13599:data <=32'h00580020;14'd13600:data <=32'h005E000E;14'd13601:data <=32'h005CFFFB;
14'd13602:data <=32'h0053FFEA;14'd13603:data <=32'h0044FFDE;14'd13604:data <=32'h0032FFD9;
14'd13605:data <=32'h0021FFDE;14'd13606:data <=32'h0014FFE8;14'd13607:data <=32'h000EFFF8;
14'd13608:data <=32'h00110009;14'd13609:data <=32'h001B0016;14'd13610:data <=32'h0029001E;
14'd13611:data <=32'h003B0022;14'd13612:data <=32'h004C001E;14'd13613:data <=32'h005E0016;
14'd13614:data <=32'h006F000A;14'd13615:data <=32'h007BFFF8;14'd13616:data <=32'h0086FFE3;
14'd13617:data <=32'h008DFFC9;14'd13618:data <=32'h008DFFAC;14'd13619:data <=32'h0085FF8D;
14'd13620:data <=32'h0076FF70;14'd13621:data <=32'h005DFF59;14'd13622:data <=32'h0040FF48;
14'd13623:data <=32'h0021FF3F;14'd13624:data <=32'h0003FF3F;14'd13625:data <=32'hFFE9FF43;
14'd13626:data <=32'hFFD5FF4A;14'd13627:data <=32'hFFC3FF50;14'd13628:data <=32'hFFB2FF54;
14'd13629:data <=32'hFF9FFF58;14'd13630:data <=32'hFF88FF5D;14'd13631:data <=32'hFF6EFF66;
14'd13632:data <=32'hFF4EFFE8;14'd13633:data <=32'hFF4DFFFA;14'd13634:data <=32'hFF4FFFFB;
14'd13635:data <=32'hFF2FFF89;14'd13636:data <=32'hFF0EFF72;14'd13637:data <=32'hFEF4FF9E;
14'd13638:data <=32'hFEE3FFCF;14'd13639:data <=32'hFEDD0004;14'd13640:data <=32'hFEE20039;
14'd13641:data <=32'hFEF2006F;14'd13642:data <=32'hFF1000A0;14'd13643:data <=32'hFF3B00CA;
14'd13644:data <=32'hFF7100E6;14'd13645:data <=32'hFFAA00F3;14'd13646:data <=32'hFFE400EC;
14'd13647:data <=32'h001500D8;14'd13648:data <=32'h003B00B7;14'd13649:data <=32'h00520091;
14'd13650:data <=32'h005B006B;14'd13651:data <=32'h005A0049;14'd13652:data <=32'h0051002E;
14'd13653:data <=32'h0042001B;14'd13654:data <=32'h0033000D;14'd13655:data <=32'h00230005;
14'd13656:data <=32'h00120003;14'd13657:data <=32'h00020006;14'd13658:data <=32'hFFF5000E;
14'd13659:data <=32'hFFEB001A;14'd13660:data <=32'hFFE90029;14'd13661:data <=32'hFFEC003A;
14'd13662:data <=32'hFFF60047;14'd13663:data <=32'h00040050;14'd13664:data <=32'h00150050;
14'd13665:data <=32'h0023004D;14'd13666:data <=32'h002D0046;14'd13667:data <=32'h0032003D;
14'd13668:data <=32'h00340036;14'd13669:data <=32'h00340032;14'd13670:data <=32'h00340032;
14'd13671:data <=32'h00370032;14'd13672:data <=32'h003F0034;14'd13673:data <=32'h00480033;
14'd13674:data <=32'h0053002E;14'd13675:data <=32'h005C0025;14'd13676:data <=32'h0063001A;
14'd13677:data <=32'h0066000C;14'd13678:data <=32'h00660001;14'd13679:data <=32'h0063FFF6;
14'd13680:data <=32'h0060FFEE;14'd13681:data <=32'h005EFFE7;14'd13682:data <=32'h005BFFE2;
14'd13683:data <=32'h0059FFDB;14'd13684:data <=32'h0056FFD5;14'd13685:data <=32'h0053FFD1;
14'd13686:data <=32'h0050FFCC;14'd13687:data <=32'h004FFFCB;14'd13688:data <=32'h0051FFC9;
14'd13689:data <=32'h0057FFC6;14'd13690:data <=32'h0061FFBE;14'd13691:data <=32'h006DFFAF;
14'd13692:data <=32'h0076FF96;14'd13693:data <=32'h0076FF75;14'd13694:data <=32'h006AFF4F;
14'd13695:data <=32'h0051FF2A;14'd13696:data <=32'hFFBFFF54;14'd13697:data <=32'hFFA8FF53;
14'd13698:data <=32'hFFA9FF5A;14'd13699:data <=32'h0000FF28;14'd13700:data <=32'hFFCDFEE8;
14'd13701:data <=32'hFF97FEF1;14'd13702:data <=32'hFF64FF05;14'd13703:data <=32'hFF36FF26;
14'd13704:data <=32'hFF0FFF4F;14'd13705:data <=32'hFEF2FF83;14'd13706:data <=32'hFEE2FFBC;
14'd13707:data <=32'hFEE2FFF9;14'd13708:data <=32'hFEF10032;14'd13709:data <=32'hFF0F0062;
14'd13710:data <=32'hFF370085;14'd13711:data <=32'hFF63009A;14'd13712:data <=32'hFF8E00A1;
14'd13713:data <=32'hFFB2009E;14'd13714:data <=32'hFFD00094;14'd13715:data <=32'hFFE70087;
14'd13716:data <=32'hFFF8007A;14'd13717:data <=32'h0006006C;14'd13718:data <=32'h0011005F;
14'd13719:data <=32'h00190050;14'd13720:data <=32'h001F0041;14'd13721:data <=32'h001F0030;
14'd13722:data <=32'h001B0022;14'd13723:data <=32'h00140017;14'd13724:data <=32'h00090011;
14'd13725:data <=32'h0000000D;14'd13726:data <=32'hFFF6000E;14'd13727:data <=32'hFFEF0012;
14'd13728:data <=32'hFFE90015;14'd13729:data <=32'hFFE30019;14'd13730:data <=32'hFFDD001E;
14'd13731:data <=32'hFFD60026;14'd13732:data <=32'hFFD00032;14'd13733:data <=32'hFFCC0042;
14'd13734:data <=32'hFFCF0057;14'd13735:data <=32'hFFD8006C;14'd13736:data <=32'hFFEA0081;
14'd13737:data <=32'h0005008F;14'd13738:data <=32'h00240094;14'd13739:data <=32'h0044008F;
14'd13740:data <=32'h00600081;14'd13741:data <=32'h0078006C;14'd13742:data <=32'h00850052;
14'd13743:data <=32'h008C0039;14'd13744:data <=32'h008D001F;14'd13745:data <=32'h0087000A;
14'd13746:data <=32'h007FFFF7;14'd13747:data <=32'h0073FFE9;14'd13748:data <=32'h0066FFDF;
14'd13749:data <=32'h0057FFDB;14'd13750:data <=32'h0049FFDB;14'd13751:data <=32'h003EFFE2;
14'd13752:data <=32'h0039FFEE;14'd13753:data <=32'h003DFFFB;14'd13754:data <=32'h004A0007;
14'd13755:data <=32'h005F000A;14'd13756:data <=32'h00790003;14'd13757:data <=32'h0091FFF0;
14'd13758:data <=32'h00A4FFD1;14'd13759:data <=32'h00ACFFAA;14'd13760:data <=32'h0087FFA8;
14'd13761:data <=32'h008DFF80;14'd13762:data <=32'h0080FF6E;14'd13763:data <=32'h0066FF8D;
14'd13764:data <=32'h004FFF40;14'd13765:data <=32'h0030FF34;14'd13766:data <=32'h0010FF2F;
14'd13767:data <=32'hFFF0FF30;14'd13768:data <=32'hFFD1FF35;14'd13769:data <=32'hFFB2FF41;
14'd13770:data <=32'hFF96FF54;14'd13771:data <=32'hFF80FF6C;14'd13772:data <=32'hFF71FF88;
14'd13773:data <=32'hFF6AFFA4;14'd13774:data <=32'hFF6BFFBC;14'd13775:data <=32'hFF6FFFCF;
14'd13776:data <=32'hFF74FFDE;14'd13777:data <=32'hFF76FFE9;14'd13778:data <=32'hFF75FFF3;
14'd13779:data <=32'hFF730000;14'd13780:data <=32'hFF720012;14'd13781:data <=32'hFF740027;
14'd13782:data <=32'hFF7D003D;14'd13783:data <=32'hFF8D0051;14'd13784:data <=32'hFFA3005F;
14'd13785:data <=32'hFFBA0067;14'd13786:data <=32'hFFD30068;14'd13787:data <=32'hFFE80063;
14'd13788:data <=32'hFFFB0058;14'd13789:data <=32'h0009004B;14'd13790:data <=32'h0014003B;
14'd13791:data <=32'h001A0029;14'd13792:data <=32'h001B0016;14'd13793:data <=32'h00150003;
14'd13794:data <=32'h0008FFF0;14'd13795:data <=32'hFFF4FFE3;14'd13796:data <=32'hFFDBFFDE;
14'd13797:data <=32'hFFC1FFE3;14'd13798:data <=32'hFFA6FFF4;14'd13799:data <=32'hFF93000C;
14'd13800:data <=32'hFF8A002D;14'd13801:data <=32'hFF8C004F;14'd13802:data <=32'hFF990070;
14'd13803:data <=32'hFFB0008A;14'd13804:data <=32'hFFCC009B;14'd13805:data <=32'hFFE900A4;
14'd13806:data <=32'h000600A5;14'd13807:data <=32'h002000A1;14'd13808:data <=32'h00370098;
14'd13809:data <=32'h004A008D;14'd13810:data <=32'h005B0080;14'd13811:data <=32'h00690071;
14'd13812:data <=32'h00740061;14'd13813:data <=32'h007A0050;14'd13814:data <=32'h007E0040;
14'd13815:data <=32'h007E0032;14'd13816:data <=32'h007D0029;14'd13817:data <=32'h007E0023;
14'd13818:data <=32'h0081001F;14'd13819:data <=32'h008A0019;14'd13820:data <=32'h0096000F;
14'd13821:data <=32'h00A3FFFE;14'd13822:data <=32'h00ACFFE6;14'd13823:data <=32'h00AEFFC9;
14'd13824:data <=32'h006F0052;14'd13825:data <=32'h00A10041;14'd13826:data <=32'h00BA0017;
14'd13827:data <=32'h0075FF9B;14'd13828:data <=32'h005AFF59;14'd13829:data <=32'h003BFF5B;
14'd13830:data <=32'h0020FF62;14'd13831:data <=32'h000CFF70;14'd13832:data <=32'hFFFDFF7D;
14'd13833:data <=32'hFFF2FF8A;14'd13834:data <=32'hFFEAFF97;14'd13835:data <=32'hFFE8FFA3;
14'd13836:data <=32'hFFE9FFB0;14'd13837:data <=32'hFFF0FFB7;14'd13838:data <=32'hFFF8FFB8;
14'd13839:data <=32'hFFFFFFB2;14'd13840:data <=32'h0002FFA5;14'd13841:data <=32'hFFFDFF96;
14'd13842:data <=32'hFFECFF85;14'd13843:data <=32'hFFD4FF7B;14'd13844:data <=32'hFFB6FF7B;
14'd13845:data <=32'hFF99FF86;14'd13846:data <=32'hFF7FFF9A;14'd13847:data <=32'hFF6EFFB6;
14'd13848:data <=32'hFF66FFD6;14'd13849:data <=32'hFF67FFF5;14'd13850:data <=32'hFF700011;
14'd13851:data <=32'hFF7E0027;14'd13852:data <=32'hFF90003A;14'd13853:data <=32'hFFA50046;
14'd13854:data <=32'hFFBC004E;14'd13855:data <=32'hFFD5004F;14'd13856:data <=32'hFFEB0048;
14'd13857:data <=32'hFFFE003B;14'd13858:data <=32'h000B0028;14'd13859:data <=32'h00110012;
14'd13860:data <=32'h000DFFFB;14'd13861:data <=32'h0001FFE9;14'd13862:data <=32'hFFEDFFDC;
14'd13863:data <=32'hFFD8FFD8;14'd13864:data <=32'hFFC2FFDC;14'd13865:data <=32'hFFAFFFE8;
14'd13866:data <=32'hFFA3FFF5;14'd13867:data <=32'hFF9B0006;14'd13868:data <=32'hFF960016;
14'd13869:data <=32'hFF950025;14'd13870:data <=32'hFF940034;14'd13871:data <=32'hFF920044;
14'd13872:data <=32'hFF920056;14'd13873:data <=32'hFF95006B;14'd13874:data <=32'hFF9C0082;
14'd13875:data <=32'hFFAA009A;14'd13876:data <=32'hFFBE00B1;14'd13877:data <=32'hFFD900C2;
14'd13878:data <=32'hFFF600D0;14'd13879:data <=32'h001700D7;14'd13880:data <=32'h003A00D9;
14'd13881:data <=32'h005D00D5;14'd13882:data <=32'h008200CD;14'd13883:data <=32'h00A700BD;
14'd13884:data <=32'h00CC00A3;14'd13885:data <=32'h00EE007E;14'd13886:data <=32'h01070051;
14'd13887:data <=32'h0113001B;14'd13888:data <=32'h002C005B;14'd13889:data <=32'h00540069;
14'd13890:data <=32'h008B0061;14'd13891:data <=32'h00EFFFDB;14'd13892:data <=32'h00D2FF7C;
14'd13893:data <=32'h00A7FF65;14'd13894:data <=32'h007CFF5C;14'd13895:data <=32'h0056FF5F;
14'd13896:data <=32'h0036FF67;14'd13897:data <=32'h001CFF74;14'd13898:data <=32'h0007FF86;
14'd13899:data <=32'hFFFAFF9A;14'd13900:data <=32'hFFF4FFB0;14'd13901:data <=32'hFFF8FFC4;
14'd13902:data <=32'h0002FFD2;14'd13903:data <=32'h0012FFD8;14'd13904:data <=32'h0022FFD4;
14'd13905:data <=32'h002DFFC7;14'd13906:data <=32'h0032FFB5;14'd13907:data <=32'h002BFFA1;
14'd13908:data <=32'h001DFF90;14'd13909:data <=32'h0007FF86;14'd13910:data <=32'hFFF0FF83;
14'd13911:data <=32'hFFDBFF89;14'd13912:data <=32'hFFC9FF94;14'd13913:data <=32'hFFBCFFA0;
14'd13914:data <=32'hFFB4FFAE;14'd13915:data <=32'hFFAEFFBB;14'd13916:data <=32'hFFAAFFC8;
14'd13917:data <=32'hFFA8FFD5;14'd13918:data <=32'hFFA8FFE2;14'd13919:data <=32'hFFAAFFEE;
14'd13920:data <=32'hFFB0FFFB;14'd13921:data <=32'hFFB90004;14'd13922:data <=32'hFFC3000A;
14'd13923:data <=32'hFFCD000B;14'd13924:data <=32'hFFD50008;14'd13925:data <=32'hFFDA0005;
14'd13926:data <=32'hFFDC0000;14'd13927:data <=32'hFFDCFFFD;14'd13928:data <=32'hFFDCFFFC;
14'd13929:data <=32'hFFDCFFFC;14'd13930:data <=32'hFFDFFFF9;14'd13931:data <=32'hFFE1FFF4;
14'd13932:data <=32'hFFE2FFEC;14'd13933:data <=32'hFFDEFFE0;14'd13934:data <=32'hFFD3FFD2;
14'd13935:data <=32'hFFC1FFC9;14'd13936:data <=32'hFFA6FFC5;14'd13937:data <=32'hFF88FFCB;
14'd13938:data <=32'hFF6BFFDB;14'd13939:data <=32'hFF50FFF7;14'd13940:data <=32'hFF3E001B;
14'd13941:data <=32'hFF350045;14'd13942:data <=32'hFF360072;14'd13943:data <=32'hFF4300A0;
14'd13944:data <=32'hFF5B00CB;14'd13945:data <=32'hFF7C00F3;14'd13946:data <=32'hFFA70114;
14'd13947:data <=32'hFFDD012C;14'd13948:data <=32'h00190139;14'd13949:data <=32'h005A0134;
14'd13950:data <=32'h009A011E;14'd13951:data <=32'h00D200F6;14'd13952:data <=32'h00450095;
14'd13953:data <=32'h0066009E;14'd13954:data <=32'h008900AC;14'd13955:data <=32'h00D300BF;
14'd13956:data <=32'h00E40058;14'd13957:data <=32'h00E00031;14'd13958:data <=32'h00D60010;
14'd13959:data <=32'h00C8FFF6;14'd13960:data <=32'h00BAFFE0;14'd13961:data <=32'h00AAFFCB;
14'd13962:data <=32'h0099FFBA;14'd13963:data <=32'h0086FFAE;14'd13964:data <=32'h0073FFA7;
14'd13965:data <=32'h0061FFA4;14'd13966:data <=32'h0054FFA5;14'd13967:data <=32'h004BFFA5;
14'd13968:data <=32'h0043FFA5;14'd13969:data <=32'h003CFFA1;14'd13970:data <=32'h0033FF9B;
14'd13971:data <=32'h0027FF95;14'd13972:data <=32'h0016FF93;14'd13973:data <=32'h0005FF95;
14'd13974:data <=32'hFFF4FF9F;14'd13975:data <=32'hFFE8FFAD;14'd13976:data <=32'hFFE3FFBD;
14'd13977:data <=32'hFFE5FFCC;14'd13978:data <=32'hFFECFFD7;14'd13979:data <=32'hFFF6FFDC;
14'd13980:data <=32'hFFFEFFDC;14'd13981:data <=32'h0005FFD7;14'd13982:data <=32'h0007FFCF;
14'd13983:data <=32'h0006FFC8;14'd13984:data <=32'h0002FFC0;14'd13985:data <=32'hFFFBFFBC;
14'd13986:data <=32'hFFF5FFB8;14'd13987:data <=32'hFFECFFB6;14'd13988:data <=32'hFFE2FFB4;
14'd13989:data <=32'hFFD6FFB6;14'd13990:data <=32'hFFCCFFBB;14'd13991:data <=32'hFFC1FFC4;
14'd13992:data <=32'hFFBAFFD1;14'd13993:data <=32'hFFB9FFE0;14'd13994:data <=32'hFFBDFFEE;
14'd13995:data <=32'hFFC8FFF7;14'd13996:data <=32'hFFD7FFFB;14'd13997:data <=32'hFFE5FFF5;
14'd13998:data <=32'hFFEEFFE7;14'd13999:data <=32'hFFF0FFD4;14'd14000:data <=32'hFFE7FFC1;
14'd14001:data <=32'hFFD4FFAF;14'd14002:data <=32'hFFBBFFA5;14'd14003:data <=32'hFF9EFFA5;
14'd14004:data <=32'hFF7FFFAF;14'd14005:data <=32'hFF63FFC1;14'd14006:data <=32'hFF4BFFDA;
14'd14007:data <=32'hFF39FFF9;14'd14008:data <=32'hFF2D001E;14'd14009:data <=32'hFF2A0046;
14'd14010:data <=32'hFF2E0070;14'd14011:data <=32'hFF3E009C;14'd14012:data <=32'hFF5900C3;
14'd14013:data <=32'hFF7E00E5;14'd14014:data <=32'hFFAB00FB;14'd14015:data <=32'hFFDC0105;
14'd14016:data <=32'hFFBE0100;14'd14017:data <=32'hFFEE011D;14'd14018:data <=32'h00100123;
14'd14019:data <=32'hFFEA00EE;14'd14020:data <=32'h000900B2;14'd14021:data <=32'h001800B2;
14'd14022:data <=32'h002900B5;14'd14023:data <=32'h003E00B7;14'd14024:data <=32'h005900B6;
14'd14025:data <=32'h007700AD;14'd14026:data <=32'h0093009C;14'd14027:data <=32'h00AD0085;
14'd14028:data <=32'h00C00068;14'd14029:data <=32'h00CE0048;14'd14030:data <=32'h00D50027;
14'd14031:data <=32'h00D80004;14'd14032:data <=32'h00D4FFE0;14'd14033:data <=32'h00C9FFBC;
14'd14034:data <=32'h00B5FF9A;14'd14035:data <=32'h0098FF7B;14'd14036:data <=32'h0073FF66;
14'd14037:data <=32'h0049FF5D;14'd14038:data <=32'h001FFF5F;14'd14039:data <=32'hFFF9FF70;
14'd14040:data <=32'hFFDDFF8C;14'd14041:data <=32'hFFCEFFAB;14'd14042:data <=32'hFFCAFFCA;
14'd14043:data <=32'hFFD1FFE6;14'd14044:data <=32'hFFE0FFFB;14'd14045:data <=32'hFFF20007;
14'd14046:data <=32'h0005000C;14'd14047:data <=32'h0017000C;14'd14048:data <=32'h00260005;
14'd14049:data <=32'h0034FFFB;14'd14050:data <=32'h003DFFEE;14'd14051:data <=32'h0043FFDE;
14'd14052:data <=32'h0044FFCC;14'd14053:data <=32'h003FFFB9;14'd14054:data <=32'h0035FFA9;
14'd14055:data <=32'h0026FF9D;14'd14056:data <=32'h0015FF96;14'd14057:data <=32'h0003FF95;
14'd14058:data <=32'hFFF5FF99;14'd14059:data <=32'hFFEBFF9F;14'd14060:data <=32'hFFE6FFA5;
14'd14061:data <=32'hFFE3FFA8;14'd14062:data <=32'hFFE2FFA7;14'd14063:data <=32'hFFDDFFA1;
14'd14064:data <=32'hFFD4FF9C;14'd14065:data <=32'hFFC5FF96;14'd14066:data <=32'hFFB3FF96;
14'd14067:data <=32'hFF9EFF9B;14'd14068:data <=32'hFF8BFFA7;14'd14069:data <=32'hFF7BFFB6;
14'd14070:data <=32'hFF70FFCA;14'd14071:data <=32'hFF69FFDE;14'd14072:data <=32'hFF66FFF2;
14'd14073:data <=32'hFF650004;14'd14074:data <=32'hFF660017;14'd14075:data <=32'hFF69002A;
14'd14076:data <=32'hFF70003C;14'd14077:data <=32'hFF7A004E;14'd14078:data <=32'hFF88005B;
14'd14079:data <=32'hFF970065;14'd14080:data <=32'hFF090081;14'd14081:data <=32'hFF1900BD;
14'd14082:data <=32'hFF4400DA;14'd14083:data <=32'hFF970060;14'd14084:data <=32'hFF99002D;
14'd14085:data <=32'hFF89003D;14'd14086:data <=32'hFF7E0057;14'd14087:data <=32'hFF7C0079;
14'd14088:data <=32'hFF87009E;14'd14089:data <=32'hFFA000BE;14'd14090:data <=32'hFFC200D9;
14'd14091:data <=32'hFFEB00EA;14'd14092:data <=32'h001700F1;14'd14093:data <=32'h004400EC;
14'd14094:data <=32'h006F00DE;14'd14095:data <=32'h009700C7;14'd14096:data <=32'h00BA00A7;
14'd14097:data <=32'h00D6007E;14'd14098:data <=32'h00E7004F;14'd14099:data <=32'h00EB001B;
14'd14100:data <=32'h00E1FFE9;14'd14101:data <=32'h00C8FFBD;14'd14102:data <=32'h00A5FF9B;
14'd14103:data <=32'h007CFF88;14'd14104:data <=32'h0054FF82;14'd14105:data <=32'h0030FF89;
14'd14106:data <=32'h0013FF98;14'd14107:data <=32'hFFFFFFAA;14'd14108:data <=32'hFFF4FFBF;
14'd14109:data <=32'hFFEEFFD2;14'd14110:data <=32'hFFEBFFE3;14'd14111:data <=32'hFFEDFFF3;
14'd14112:data <=32'hFFF30003;14'd14113:data <=32'hFFFC0010;14'd14114:data <=32'h0008001A;
14'd14115:data <=32'h00180022;14'd14116:data <=32'h002B0024;14'd14117:data <=32'h003D0020;
14'd14118:data <=32'h004D0016;14'd14119:data <=32'h005B0009;14'd14120:data <=32'h0066FFF9;
14'd14121:data <=32'h006DFFE7;14'd14122:data <=32'h0070FFD5;14'd14123:data <=32'h0073FFC1;
14'd14124:data <=32'h0072FFAC;14'd14125:data <=32'h006EFF95;14'd14126:data <=32'h0066FF7A;
14'd14127:data <=32'h0056FF5F;14'd14128:data <=32'h003DFF46;14'd14129:data <=32'h001AFF32;
14'd14130:data <=32'hFFF2FF28;14'd14131:data <=32'hFFC5FF29;14'd14132:data <=32'hFF9BFF37;
14'd14133:data <=32'hFF76FF50;14'd14134:data <=32'hFF5BFF71;14'd14135:data <=32'hFF4AFF96;
14'd14136:data <=32'hFF44FFBB;14'd14137:data <=32'hFF46FFDD;14'd14138:data <=32'hFF4EFFFA;
14'd14139:data <=32'hFF5D0014;14'd14140:data <=32'hFF6E0028;14'd14141:data <=32'hFF830036;
14'd14142:data <=32'hFF99003C;14'd14143:data <=32'hFFAE003C;14'd14144:data <=32'hFF47FFD1;
14'd14145:data <=32'hFF30FFEF;14'd14146:data <=32'hFF34001D;14'd14147:data <=32'hFFA5003F;
14'd14148:data <=32'hFFAEFFFB;14'd14149:data <=32'hFF9BFFF9;14'd14150:data <=32'hFF870002;
14'd14151:data <=32'hFF750015;14'd14152:data <=32'hFF6A0031;14'd14153:data <=32'hFF69004F;
14'd14154:data <=32'hFF73006E;14'd14155:data <=32'hFF83008A;14'd14156:data <=32'hFF9A009E;
14'd14157:data <=32'hFFB400AF;14'd14158:data <=32'hFFD000BA;14'd14159:data <=32'hFFEF00C0;
14'd14160:data <=32'h000F00C1;14'd14161:data <=32'h003000BA;14'd14162:data <=32'h004F00AC;
14'd14163:data <=32'h00690095;14'd14164:data <=32'h007D0079;14'd14165:data <=32'h0085005A;
14'd14166:data <=32'h0086003C;14'd14167:data <=32'h007F0024;14'd14168:data <=32'h00750011;
14'd14169:data <=32'h00690005;14'd14170:data <=32'h005FFFFD;14'd14171:data <=32'h0057FFF6;
14'd14172:data <=32'h0051FFEF;14'd14173:data <=32'h004AFFE7;14'd14174:data <=32'h0040FFDE;
14'd14175:data <=32'h0033FFD8;14'd14176:data <=32'h0023FFD6;14'd14177:data <=32'h0013FFDA;
14'd14178:data <=32'h0003FFE4;14'd14179:data <=32'hFFF9FFF2;14'd14180:data <=32'hFFF40004;
14'd14181:data <=32'hFFF50017;14'd14182:data <=32'hFFFD0028;14'd14183:data <=32'h000B0038;
14'd14184:data <=32'h001D0044;14'd14185:data <=32'h0033004B;14'd14186:data <=32'h004C004E;
14'd14187:data <=32'h0069004B;14'd14188:data <=32'h0086003E;14'd14189:data <=32'h00A30029;
14'd14190:data <=32'h00BB000A;14'd14191:data <=32'h00CCFFE0;14'd14192:data <=32'h00D0FFAF;
14'd14193:data <=32'h00C6FF7D;14'd14194:data <=32'h00ADFF4F;14'd14195:data <=32'h0086FF29;
14'd14196:data <=32'h0057FF10;14'd14197:data <=32'h0026FF04;14'd14198:data <=32'hFFF5FF09;
14'd14199:data <=32'hFFC9FF15;14'd14200:data <=32'hFFA5FF2B;14'd14201:data <=32'hFF88FF45;
14'd14202:data <=32'hFF73FF61;14'd14203:data <=32'hFF66FF7F;14'd14204:data <=32'hFF5EFF9D;
14'd14205:data <=32'hFF5DFFBA;14'd14206:data <=32'hFF63FFD5;14'd14207:data <=32'hFF6EFFEA;
14'd14208:data <=32'hFF9DFFD7;14'd14209:data <=32'hFF99FFD6;14'd14210:data <=32'hFF86FFDE;
14'd14211:data <=32'hFF53FFF5;14'd14212:data <=32'hFF61FFC9;14'd14213:data <=32'hFF56FFDA;
14'd14214:data <=32'hFF4CFFEE;14'd14215:data <=32'hFF460009;14'd14216:data <=32'hFF470028;
14'd14217:data <=32'hFF510048;14'd14218:data <=32'hFF640062;14'd14219:data <=32'hFF7E0076;
14'd14220:data <=32'hFF990081;14'd14221:data <=32'hFFB30085;14'd14222:data <=32'hFFCA0082;
14'd14223:data <=32'hFFDC007E;14'd14224:data <=32'hFFEC0076;14'd14225:data <=32'hFFF9006E;
14'd14226:data <=32'h00040065;14'd14227:data <=32'h000B005B;14'd14228:data <=32'h000F004F;
14'd14229:data <=32'h000F0045;14'd14230:data <=32'h000C003D;14'd14231:data <=32'h0006003B;
14'd14232:data <=32'h0000003E;14'd14233:data <=32'hFFFF0046;14'd14234:data <=32'h00040051;
14'd14235:data <=32'h00100059;14'd14236:data <=32'h001F005B;14'd14237:data <=32'h00320059;
14'd14238:data <=32'h0042004D;14'd14239:data <=32'h004E003B;14'd14240:data <=32'h00500027;
14'd14241:data <=32'h004D0014;14'd14242:data <=32'h00420006;14'd14243:data <=32'h0035FFFC;
14'd14244:data <=32'h0026FFF9;14'd14245:data <=32'h0018FFFB;14'd14246:data <=32'h000C0002;
14'd14247:data <=32'h0002000C;14'd14248:data <=32'hFFFE001B;14'd14249:data <=32'hFFFE002B;
14'd14250:data <=32'h0004003D;14'd14251:data <=32'h000F004F;14'd14252:data <=32'h0023005D;
14'd14253:data <=32'h003D0066;14'd14254:data <=32'h005B0067;14'd14255:data <=32'h007C005D;
14'd14256:data <=32'h009A0049;14'd14257:data <=32'h00B1002C;14'd14258:data <=32'h00BF0008;
14'd14259:data <=32'h00C1FFE3;14'd14260:data <=32'h00BBFFC1;14'd14261:data <=32'h00ADFFA3;
14'd14262:data <=32'h009DFF8C;14'd14263:data <=32'h008AFF79;14'd14264:data <=32'h0078FF69;
14'd14265:data <=32'h0067FF5C;14'd14266:data <=32'h0053FF4E;14'd14267:data <=32'h003EFF41;
14'd14268:data <=32'h0026FF37;14'd14269:data <=32'h000BFF30;14'd14270:data <=32'hFFEFFF2F;
14'd14271:data <=32'hFFD3FF33;14'd14272:data <=32'hFF91FFAE;14'd14273:data <=32'hFF97FFB9;
14'd14274:data <=32'hFFA1FFAD;14'd14275:data <=32'hFF9EFF30;14'd14276:data <=32'hFF87FF01;
14'd14277:data <=32'hFF57FF17;14'd14278:data <=32'hFF2BFF39;14'd14279:data <=32'hFF06FF66;
14'd14280:data <=32'hFEF0FF9E;14'd14281:data <=32'hFEE9FFDB;14'd14282:data <=32'hFEF40015;
14'd14283:data <=32'hFF0E0048;14'd14284:data <=32'hFF31006E;14'd14285:data <=32'hFF5B0087;
14'd14286:data <=32'hFF850093;14'd14287:data <=32'hFFAC0094;14'd14288:data <=32'hFFCE008D;
14'd14289:data <=32'hFFEA007F;14'd14290:data <=32'h0001006D;14'd14291:data <=32'h00100056;
14'd14292:data <=32'h00180040;14'd14293:data <=32'h00170028;14'd14294:data <=32'h000D0012;
14'd14295:data <=32'hFFFD0006;14'd14296:data <=32'hFFEA0001;14'd14297:data <=32'hFFD70006;
14'd14298:data <=32'hFFC80013;14'd14299:data <=32'hFFC30026;14'd14300:data <=32'hFFC50038;
14'd14301:data <=32'hFFCE0047;14'd14302:data <=32'hFFDC0052;14'd14303:data <=32'hFFEA0055;
14'd14304:data <=32'hFFF70053;14'd14305:data <=32'h00010050;14'd14306:data <=32'h0007004A;
14'd14307:data <=32'h000B0046;14'd14308:data <=32'h000E0044;14'd14309:data <=32'h00100043;
14'd14310:data <=32'h00130042;14'd14311:data <=32'h00170040;14'd14312:data <=32'h0019003F;
14'd14313:data <=32'h001C003D;14'd14314:data <=32'h001E003D;14'd14315:data <=32'h001F003E;
14'd14316:data <=32'h00220042;14'd14317:data <=32'h00280045;14'd14318:data <=32'h00300048;
14'd14319:data <=32'h003C0047;14'd14320:data <=32'h00460044;14'd14321:data <=32'h0051003D;
14'd14322:data <=32'h00560035;14'd14323:data <=32'h005A002B;14'd14324:data <=32'h005A0026;
14'd14325:data <=32'h005B0024;14'd14326:data <=32'h005F0026;14'd14327:data <=32'h00690029;
14'd14328:data <=32'h0078002A;14'd14329:data <=32'h008E0024;14'd14330:data <=32'h00A60015;
14'd14331:data <=32'h00BBFFFC;14'd14332:data <=32'h00CBFFDB;14'd14333:data <=32'h00D2FFB4;
14'd14334:data <=32'h00CFFF8A;14'd14335:data <=32'h00C3FF60;14'd14336:data <=32'h0017FF65;
14'd14337:data <=32'h0011FF61;14'd14338:data <=32'h0020FF65;14'd14339:data <=32'h0090FF3D;
14'd14340:data <=32'h007BFEE2;14'd14341:data <=32'h0041FEC8;14'd14342:data <=32'hFFFFFEBF;
14'd14343:data <=32'hFFBCFEC6;14'd14344:data <=32'hFF7EFEE0;14'd14345:data <=32'hFF4BFF0A;
14'd14346:data <=32'hFF27FF3F;14'd14347:data <=32'hFF14FF77;14'd14348:data <=32'hFF11FFAD;
14'd14349:data <=32'hFF1BFFDC;14'd14350:data <=32'hFF2B0003;14'd14351:data <=32'hFF410022;
14'd14352:data <=32'hFF5A003A;14'd14353:data <=32'hFF73004B;14'd14354:data <=32'hFF8F0057;
14'd14355:data <=32'hFFAA005B;14'd14356:data <=32'hFFC40058;14'd14357:data <=32'hFFDA004F;
14'd14358:data <=32'hFFEA0041;14'd14359:data <=32'hFFF20031;14'd14360:data <=32'hFFF50023;
14'd14361:data <=32'hFFF10018;14'd14362:data <=32'hFFEB0012;14'd14363:data <=32'hFFE50010;
14'd14364:data <=32'hFFE30010;14'd14365:data <=32'hFFE10010;14'd14366:data <=32'hFFE1000F;
14'd14367:data <=32'hFFE0000C;14'd14368:data <=32'hFFDB0007;14'd14369:data <=32'hFFD30005;
14'd14370:data <=32'hFFC70006;14'd14371:data <=32'hFFBB000D;14'd14372:data <=32'hFFB0001B;
14'd14373:data <=32'hFFAA002C;14'd14374:data <=32'hFFAA0041;14'd14375:data <=32'hFFB10056;
14'd14376:data <=32'hFFBD0067;14'd14377:data <=32'hFFCE0074;14'd14378:data <=32'hFFE1007E;
14'd14379:data <=32'hFFF50082;14'd14380:data <=32'h00090081;14'd14381:data <=32'h001C007E;
14'd14382:data <=32'h002E0077;14'd14383:data <=32'h003F006B;14'd14384:data <=32'h004B005C;
14'd14385:data <=32'h0052004A;14'd14386:data <=32'h00530036;14'd14387:data <=32'h004A0026;
14'd14388:data <=32'h003E001B;14'd14389:data <=32'h002E001A;14'd14390:data <=32'h00200023;
14'd14391:data <=32'h00180034;14'd14392:data <=32'h001C0048;14'd14393:data <=32'h002A005D;
14'd14394:data <=32'h0044006D;14'd14395:data <=32'h00640072;14'd14396:data <=32'h0087006D;
14'd14397:data <=32'h00AA005C;14'd14398:data <=32'h00C70041;14'd14399:data <=32'h00DF001F;
14'd14400:data <=32'h00A50000;14'd14401:data <=32'h00BFFFE8;14'd14402:data <=32'h00C9FFDB;
14'd14403:data <=32'h00C2FFF3;14'd14404:data <=32'h00D6FF95;14'd14405:data <=32'h00C1FF6D;
14'd14406:data <=32'h00A3FF4C;14'd14407:data <=32'h007FFF33;14'd14408:data <=32'h0055FF26;
14'd14409:data <=32'h002AFF24;14'd14410:data <=32'h0006FF2D;14'd14411:data <=32'hFFEAFF3B;
14'd14412:data <=32'hFFD5FF4B;14'd14413:data <=32'hFFC5FF5A;14'd14414:data <=32'hFFB8FF68;
14'd14415:data <=32'hFFABFF74;14'd14416:data <=32'hFF9DFF80;14'd14417:data <=32'hFF8FFF8F;
14'd14418:data <=32'hFF83FFA2;14'd14419:data <=32'hFF7BFFB7;14'd14420:data <=32'hFF78FFCD;
14'd14421:data <=32'hFF79FFE3;14'd14422:data <=32'hFF7EFFF6;14'd14423:data <=32'hFF860007;
14'd14424:data <=32'hFF900016;14'd14425:data <=32'hFF9A0024;14'd14426:data <=32'hFFA7002F;
14'd14427:data <=32'hFFBA003A;14'd14428:data <=32'hFFCC003F;14'd14429:data <=32'hFFE2003E;
14'd14430:data <=32'hFFF80035;14'd14431:data <=32'h000A0025;14'd14432:data <=32'h0013000E;
14'd14433:data <=32'h0013FFF4;14'd14434:data <=32'h0007FFDC;14'd14435:data <=32'hFFF3FFCA;
14'd14436:data <=32'hFFD9FFC1;14'd14437:data <=32'hFFBDFFC2;14'd14438:data <=32'hFFA3FFCE;
14'd14439:data <=32'hFF8EFFE1;14'd14440:data <=32'hFF7FFFF9;14'd14441:data <=32'hFF790013;
14'd14442:data <=32'hFF78002D;14'd14443:data <=32'hFF7D0047;14'd14444:data <=32'hFF89005F;
14'd14445:data <=32'hFF980073;14'd14446:data <=32'hFFAD0085;14'd14447:data <=32'hFFC50091;
14'd14448:data <=32'hFFDE0095;14'd14449:data <=32'hFFF70093;14'd14450:data <=32'h000C0089;
14'd14451:data <=32'h001B007D;14'd14452:data <=32'h00220070;14'd14453:data <=32'h00230064;
14'd14454:data <=32'h00220060;14'd14455:data <=32'h001F0063;14'd14456:data <=32'h0021006A;
14'd14457:data <=32'h00290074;14'd14458:data <=32'h0039007C;14'd14459:data <=32'h004E007E;
14'd14460:data <=32'h0066007B;14'd14461:data <=32'h007C0070;14'd14462:data <=32'h00910060;
14'd14463:data <=32'h00A1004C;14'd14464:data <=32'h003800A2;14'd14465:data <=32'h007000B1;
14'd14466:data <=32'h009D009E;14'd14467:data <=32'h008F0022;14'd14468:data <=32'h00A4FFD8;
14'd14469:data <=32'h0095FFC4;14'd14470:data <=32'h0082FFB6;14'd14471:data <=32'h006FFFAC;
14'd14472:data <=32'h005BFFA9;14'd14473:data <=32'h004AFFAD;14'd14474:data <=32'h0040FFB6;
14'd14475:data <=32'h003DFFC0;14'd14476:data <=32'h0042FFC5;14'd14477:data <=32'h004CFFC2;
14'd14478:data <=32'h0055FFB7;14'd14479:data <=32'h0058FFA6;14'd14480:data <=32'h0054FF8E;
14'd14481:data <=32'h0047FF79;14'd14482:data <=32'h0031FF67;14'd14483:data <=32'h0017FF5B;
14'd14484:data <=32'hFFFAFF57;14'd14485:data <=32'hFFDDFF5A;14'd14486:data <=32'hFFC2FF65;
14'd14487:data <=32'hFFA8FF73;14'd14488:data <=32'hFF92FF87;14'd14489:data <=32'hFF81FFA1;
14'd14490:data <=32'hFF76FFBF;14'd14491:data <=32'hFF74FFDF;14'd14492:data <=32'hFF7BFFFF;
14'd14493:data <=32'hFF8D001C;14'd14494:data <=32'hFFA7002F;14'd14495:data <=32'hFFC60038;
14'd14496:data <=32'hFFE40037;14'd14497:data <=32'hFFFD002A;14'd14498:data <=32'h000E0015;
14'd14499:data <=32'h0016FFFD;14'd14500:data <=32'h0013FFE6;14'd14501:data <=32'h0009FFD4;
14'd14502:data <=32'hFFFCFFC6;14'd14503:data <=32'hFFECFFBD;14'd14504:data <=32'hFFDAFFB8;
14'd14505:data <=32'hFFC8FFB8;14'd14506:data <=32'hFFB7FFBB;14'd14507:data <=32'hFFA6FFBF;
14'd14508:data <=32'hFF94FFC8;14'd14509:data <=32'hFF84FFD5;14'd14510:data <=32'hFF75FFE7;
14'd14511:data <=32'hFF6BFFFC;14'd14512:data <=32'hFF650013;14'd14513:data <=32'hFF64002B;
14'd14514:data <=32'hFF660042;14'd14515:data <=32'hFF6C0057;14'd14516:data <=32'hFF73006D;
14'd14517:data <=32'hFF7B0081;14'd14518:data <=32'hFF870099;14'd14519:data <=32'hFF9700B2;
14'd14520:data <=32'hFFAD00CB;14'd14521:data <=32'hFFCC00E1;14'd14522:data <=32'hFFF400F1;
14'd14523:data <=32'h002200F7;14'd14524:data <=32'h005200EF;14'd14525:data <=32'h007D00DA;
14'd14526:data <=32'h00A200BA;14'd14527:data <=32'h00BB0095;14'd14528:data <=32'hFFCE007A;
14'd14529:data <=32'hFFE800A8;14'd14530:data <=32'h002100C3;14'd14531:data <=32'h00B6006A;
14'd14532:data <=32'h00CE000F;14'd14533:data <=32'h00BCFFED;14'd14534:data <=32'h00A2FFD2;
14'd14535:data <=32'h0085FFC0;14'd14536:data <=32'h0066FFB9;14'd14537:data <=32'h0049FFBD;
14'd14538:data <=32'h0033FFCB;14'd14539:data <=32'h0027FFDF;14'd14540:data <=32'h0028FFF4;
14'd14541:data <=32'h00330004;14'd14542:data <=32'h0045000A;14'd14543:data <=32'h00590005;
14'd14544:data <=32'h006AFFF8;14'd14545:data <=32'h0074FFE3;14'd14546:data <=32'h0075FFCC;
14'd14547:data <=32'h0070FFB5;14'd14548:data <=32'h0066FFA1;14'd14549:data <=32'h0056FF90;
14'd14550:data <=32'h0045FF83;14'd14551:data <=32'h0030FF79;14'd14552:data <=32'h0019FF73;
14'd14553:data <=32'h0001FF72;14'd14554:data <=32'hFFE9FF79;14'd14555:data <=32'hFFD2FF85;
14'd14556:data <=32'hFFC1FF97;14'd14557:data <=32'hFFB6FFAE;14'd14558:data <=32'hFFB4FFC5;
14'd14559:data <=32'hFFB8FFD8;14'd14560:data <=32'hFFC2FFE6;14'd14561:data <=32'hFFCEFFF0;
14'd14562:data <=32'hFFD8FFF2;14'd14563:data <=32'hFFE1FFF2;14'd14564:data <=32'hFFE6FFF0;
14'd14565:data <=32'hFFE9FFEF;14'd14566:data <=32'hFFEDFFEF;14'd14567:data <=32'hFFF2FFEF;
14'd14568:data <=32'hFFF8FFED;14'd14569:data <=32'h0000FFE7;14'd14570:data <=32'h0007FFDE;
14'd14571:data <=32'h000BFFCF;14'd14572:data <=32'h0009FFBC;14'd14573:data <=32'h0001FFAA;
14'd14574:data <=32'hFFF0FF99;14'd14575:data <=32'hFFDAFF8B;14'd14576:data <=32'hFFBEFF84;
14'd14577:data <=32'hFFA0FF82;14'd14578:data <=32'hFF80FF88;14'd14579:data <=32'hFF60FF95;
14'd14580:data <=32'hFF40FFA9;14'd14581:data <=32'hFF22FFC7;14'd14582:data <=32'hFF08FFEE;
14'd14583:data <=32'hFEF7001F;14'd14584:data <=32'hFEF10057;14'd14585:data <=32'hFEFC0093;
14'd14586:data <=32'hFF1800CD;14'd14587:data <=32'hFF4500FF;14'd14588:data <=32'hFF7E0121;
14'd14589:data <=32'hFFBD0134;14'd14590:data <=32'hFFFD0134;14'd14591:data <=32'h00380124;
14'd14592:data <=32'hFFD20084;14'd14593:data <=32'hFFDC00A2;14'd14594:data <=32'hFFEF00CE;
14'd14595:data <=32'h0042010C;14'd14596:data <=32'h008200BD;14'd14597:data <=32'h0094009B;
14'd14598:data <=32'h009D0079;14'd14599:data <=32'h009F0059;14'd14600:data <=32'h0099003C;
14'd14601:data <=32'h008D0026;14'd14602:data <=32'h007F0018;14'd14603:data <=32'h00730011;
14'd14604:data <=32'h006B000F;14'd14605:data <=32'h0069000F;14'd14606:data <=32'h006D000C;
14'd14607:data <=32'h00720004;14'd14608:data <=32'h0075FFF7;14'd14609:data <=32'h0073FFE7;
14'd14610:data <=32'h006BFFD7;14'd14611:data <=32'h0060FFCC;14'd14612:data <=32'h0053FFC4;
14'd14613:data <=32'h0046FFC1;14'd14614:data <=32'h003BFFC1;14'd14615:data <=32'h0034FFC4;
14'd14616:data <=32'h002DFFC5;14'd14617:data <=32'h002AFFC6;14'd14618:data <=32'h0024FFC6;
14'd14619:data <=32'h0020FFC8;14'd14620:data <=32'h001BFFC9;14'd14621:data <=32'h001AFFCC;
14'd14622:data <=32'h001BFFCE;14'd14623:data <=32'h001CFFCE;14'd14624:data <=32'h001EFFCB;
14'd14625:data <=32'h001FFFC5;14'd14626:data <=32'h001CFFBB;14'd14627:data <=32'h0014FFB4;
14'd14628:data <=32'h0008FFAF;14'd14629:data <=32'hFFF9FFAF;14'd14630:data <=32'hFFEBFFB5;
14'd14631:data <=32'hFFE1FFC1;14'd14632:data <=32'hFFDEFFD1;14'd14633:data <=32'hFFE2FFDF;
14'd14634:data <=32'hFFEDFFEA;14'd14635:data <=32'hFFFDFFEE;14'd14636:data <=32'h000DFFEA;
14'd14637:data <=32'h001AFFDE;14'd14638:data <=32'h0023FFCD;14'd14639:data <=32'h0025FFB7;
14'd14640:data <=32'h0021FFA2;14'd14641:data <=32'h0014FF8A;14'd14642:data <=32'h0002FF75;
14'd14643:data <=32'hFFE9FF64;14'd14644:data <=32'hFFC9FF57;14'd14645:data <=32'hFFA1FF52;
14'd14646:data <=32'hFF77FF57;14'd14647:data <=32'hFF4BFF69;14'd14648:data <=32'hFF23FF89;
14'd14649:data <=32'hFF03FFB6;14'd14650:data <=32'hFEF1FFEA;14'd14651:data <=32'hFEED0022;
14'd14652:data <=32'hFEF90057;14'd14653:data <=32'hFF120087;14'd14654:data <=32'hFF3400AA;
14'd14655:data <=32'hFF5900C4;14'd14656:data <=32'hFF5200A3;14'd14657:data <=32'hFF6400CB;
14'd14658:data <=32'hFF6F00E6;14'd14659:data <=32'hFF5500C6;14'd14660:data <=32'hFF8E00A7;
14'd14661:data <=32'hFFA300B5;14'd14662:data <=32'hFFBB00C1;14'd14663:data <=32'hFFD600C9;
14'd14664:data <=32'hFFF000CD;14'd14665:data <=32'h000A00CC;14'd14666:data <=32'h002300CB;
14'd14667:data <=32'h003E00C7;14'd14668:data <=32'h005B00BF;14'd14669:data <=32'h007900B2;
14'd14670:data <=32'h0097009D;14'd14671:data <=32'h00B2007F;14'd14672:data <=32'h00C40059;
14'd14673:data <=32'h00CB002C;14'd14674:data <=32'h00C50001;14'd14675:data <=32'h00B3FFDB;
14'd14676:data <=32'h0097FFBD;14'd14677:data <=32'h0077FFAB;14'd14678:data <=32'h0055FFA5;
14'd14679:data <=32'h0038FFA8;14'd14680:data <=32'h0020FFB1;14'd14681:data <=32'h000DFFBF;
14'd14682:data <=32'h0001FFCF;14'd14683:data <=32'hFFFAFFE1;14'd14684:data <=32'hFFF9FFF5;
14'd14685:data <=32'hFFFE0005;14'd14686:data <=32'h000A0014;14'd14687:data <=32'h0019001D;
14'd14688:data <=32'h002E0020;14'd14689:data <=32'h0041001B;14'd14690:data <=32'h0052000D;
14'd14691:data <=32'h005CFFFB;14'd14692:data <=32'h005EFFE5;14'd14693:data <=32'h0059FFD2;
14'd14694:data <=32'h004DFFC4;14'd14695:data <=32'h0040FFBB;14'd14696:data <=32'h0033FFB8;
14'd14697:data <=32'h002AFFBA;14'd14698:data <=32'h0024FFBE;14'd14699:data <=32'h0025FFC0;
14'd14700:data <=32'h0026FFBF;14'd14701:data <=32'h0027FFBA;14'd14702:data <=32'h0028FFB2;
14'd14703:data <=32'h0025FFA9;14'd14704:data <=32'h0020FF9F;14'd14705:data <=32'h0018FF95;
14'd14706:data <=32'h000FFF8C;14'd14707:data <=32'h0004FF84;14'd14708:data <=32'hFFF6FF7C;
14'd14709:data <=32'hFFE5FF75;14'd14710:data <=32'hFFD0FF72;14'd14711:data <=32'hFFB8FF71;
14'd14712:data <=32'hFF9FFF78;14'd14713:data <=32'hFF87FF87;14'd14714:data <=32'hFF74FF9B;
14'd14715:data <=32'hFF69FFB2;14'd14716:data <=32'hFF64FFCA;14'd14717:data <=32'hFF65FFDF;
14'd14718:data <=32'hFF69FFED;14'd14719:data <=32'hFF6CFFF8;14'd14720:data <=32'hFEEFFFEE;
14'd14721:data <=32'hFEDE0022;14'd14722:data <=32'hFEEB0048;14'd14723:data <=32'hFF4DFFF7;
14'd14724:data <=32'hFF5EFFD6;14'd14725:data <=32'hFF49FFEC;14'd14726:data <=32'hFF390008;
14'd14727:data <=32'hFF30002D;14'd14728:data <=32'hFF2F0052;14'd14729:data <=32'hFF360079;
14'd14730:data <=32'hFF4500A0;14'd14731:data <=32'hFF5E00C7;14'd14732:data <=32'hFF8300E9;
14'd14733:data <=32'hFFAF0102;14'd14734:data <=32'hFFE70111;14'd14735:data <=32'h00200110;
14'd14736:data <=32'h005800FE;14'd14737:data <=32'h008800DC;14'd14738:data <=32'h00AB00B0;
14'd14739:data <=32'h00BE007E;14'd14740:data <=32'h00C2004B;14'd14741:data <=32'h00B90020;
14'd14742:data <=32'h00A6FFFC;14'd14743:data <=32'h008EFFE0;14'd14744:data <=32'h0074FFCE;
14'd14745:data <=32'h0059FFC3;14'd14746:data <=32'h003EFFBF;14'd14747:data <=32'h0025FFC1;
14'd14748:data <=32'h000EFFCA;14'd14749:data <=32'hFFFBFFD9;14'd14750:data <=32'hFFEFFFED;
14'd14751:data <=32'hFFEB0002;14'd14752:data <=32'hFFEE0018;14'd14753:data <=32'hFFF80029;
14'd14754:data <=32'h00070035;14'd14755:data <=32'h0019003B;14'd14756:data <=32'h0028003C;
14'd14757:data <=32'h00360039;14'd14758:data <=32'h00420035;14'd14759:data <=32'h004C0030;
14'd14760:data <=32'h0058002B;14'd14761:data <=32'h00650025;14'd14762:data <=32'h0074001D;
14'd14763:data <=32'h0083000F;14'd14764:data <=32'h0091FFFA;14'd14765:data <=32'h009BFFDF;
14'd14766:data <=32'h009DFFC1;14'd14767:data <=32'h0096FFA1;14'd14768:data <=32'h0087FF84;
14'd14769:data <=32'h0071FF6A;14'd14770:data <=32'h0056FF58;14'd14771:data <=32'h0038FF4D;
14'd14772:data <=32'h001AFF47;14'd14773:data <=32'hFFFCFF49;14'd14774:data <=32'hFFDFFF4E;
14'd14775:data <=32'hFFC5FF5B;14'd14776:data <=32'hFFAEFF6D;14'd14777:data <=32'hFF9CFF83;
14'd14778:data <=32'hFF92FF9D;14'd14779:data <=32'hFF91FFB8;14'd14780:data <=32'hFF9AFFCF;
14'd14781:data <=32'hFFA9FFDE;14'd14782:data <=32'hFFBBFFE4;14'd14783:data <=32'hFFCBFFDD;
14'd14784:data <=32'hFF84FF5F;14'd14785:data <=32'hFF5DFF66;14'd14786:data <=32'hFF47FF8A;
14'd14787:data <=32'hFFA3FFCC;14'd14788:data <=32'hFFB9FF96;14'd14789:data <=32'hFFA0FF94;
14'd14790:data <=32'hFF84FF98;14'd14791:data <=32'hFF6AFFA8;14'd14792:data <=32'hFF53FFBC;
14'd14793:data <=32'hFF3FFFD6;14'd14794:data <=32'hFF31FFF5;14'd14795:data <=32'hFF29001B;
14'd14796:data <=32'hFF2A0043;14'd14797:data <=32'hFF35006D;14'd14798:data <=32'hFF4D0095;
14'd14799:data <=32'hFF7000B4;14'd14800:data <=32'hFF9A00C8;14'd14801:data <=32'hFFC600CF;
14'd14802:data <=32'hFFEE00C9;14'd14803:data <=32'h001100B9;14'd14804:data <=32'h002B00A5;
14'd14805:data <=32'h003D008F;14'd14806:data <=32'h0048007B;14'd14807:data <=32'h00500067;
14'd14808:data <=32'h00550056;14'd14809:data <=32'h005A0044;14'd14810:data <=32'h005A0032;
14'd14811:data <=32'h00580020;14'd14812:data <=32'h0051000F;14'd14813:data <=32'h00460000;
14'd14814:data <=32'h0037FFF5;14'd14815:data <=32'h0028FFF1;14'd14816:data <=32'h0019FFF2;
14'd14817:data <=32'h000BFFF5;14'd14818:data <=32'h0000FFFC;14'd14819:data <=32'hFFF70004;
14'd14820:data <=32'hFFEF000E;14'd14821:data <=32'hFFE9001C;14'd14822:data <=32'hFFE5002C;
14'd14823:data <=32'hFFE60041;14'd14824:data <=32'hFFEE0057;14'd14825:data <=32'hFFFE006E;
14'd14826:data <=32'h00180082;14'd14827:data <=32'h003B008D;14'd14828:data <=32'h0062008E;
14'd14829:data <=32'h008C0081;14'd14830:data <=32'h00B20068;14'd14831:data <=32'h00CF0043;
14'd14832:data <=32'h00E00018;14'd14833:data <=32'h00E5FFEB;14'd14834:data <=32'h00DFFFBE;
14'd14835:data <=32'h00CFFF95;14'd14836:data <=32'h00B7FF71;14'd14837:data <=32'h0099FF54;
14'd14838:data <=32'h0075FF41;14'd14839:data <=32'h0050FF33;14'd14840:data <=32'h0028FF30;
14'd14841:data <=32'h0002FF37;14'd14842:data <=32'hFFE2FF47;14'd14843:data <=32'hFFC8FF5E;
14'd14844:data <=32'hFFBAFF79;14'd14845:data <=32'hFFB8FF93;14'd14846:data <=32'hFFBEFFA7;
14'd14847:data <=32'hFFC9FFB2;14'd14848:data <=32'hFFF6FFA5;14'd14849:data <=32'hFFF4FF92;
14'd14850:data <=32'hFFDBFF88;14'd14851:data <=32'hFF9CFF94;14'd14852:data <=32'hFFB3FF6D;
14'd14853:data <=32'hFF9DFF76;14'd14854:data <=32'hFF88FF84;14'd14855:data <=32'hFF77FF98;
14'd14856:data <=32'hFF6DFFAD;14'd14857:data <=32'hFF66FFC2;14'd14858:data <=32'hFF61FFD8;
14'd14859:data <=32'hFF60FFED;14'd14860:data <=32'hFF620002;14'd14861:data <=32'hFF670019;
14'd14862:data <=32'hFF73002E;14'd14863:data <=32'hFF830040;14'd14864:data <=32'hFF96004B;
14'd14865:data <=32'hFFAA004E;14'd14866:data <=32'hFFBB004D;14'd14867:data <=32'hFFC70046;
14'd14868:data <=32'hFFCB003F;14'd14869:data <=32'hFFCB003A;14'd14870:data <=32'hFFC7003B;
14'd14871:data <=32'hFFC50042;14'd14872:data <=32'hFFC7004D;14'd14873:data <=32'hFFCE0059;
14'd14874:data <=32'hFFDB0062;14'd14875:data <=32'hFFEB0067;14'd14876:data <=32'hFFFD0067;
14'd14877:data <=32'h000E0061;14'd14878:data <=32'h001C0057;14'd14879:data <=32'h0025004B;
14'd14880:data <=32'h002B003E;14'd14881:data <=32'h002E002F;14'd14882:data <=32'h002D0020;
14'd14883:data <=32'h00270012;14'd14884:data <=32'h001D0006;14'd14885:data <=32'h000EFFFE;
14'd14886:data <=32'hFFF9FFFB;14'd14887:data <=32'hFFE50002;14'd14888:data <=32'hFFD20012;
14'd14889:data <=32'hFFC60029;14'd14890:data <=32'hFFC20047;14'd14891:data <=32'hFFCB0067;
14'd14892:data <=32'hFFDF0082;14'd14893:data <=32'hFFFC0097;14'd14894:data <=32'h001F00A2;
14'd14895:data <=32'h004400A2;14'd14896:data <=32'h00660098;14'd14897:data <=32'h00830087;
14'd14898:data <=32'h009C0071;14'd14899:data <=32'h00AE0057;14'd14900:data <=32'h00BD003C;
14'd14901:data <=32'h00C7001F;14'd14902:data <=32'h00CB0001;14'd14903:data <=32'h00CBFFE2;
14'd14904:data <=32'h00C3FFC4;14'd14905:data <=32'h00B7FFA9;14'd14906:data <=32'h00A6FF92;
14'd14907:data <=32'h0093FF81;14'd14908:data <=32'h0080FF74;14'd14909:data <=32'h0070FF6B;
14'd14910:data <=32'h0062FF61;14'd14911:data <=32'h0054FF55;14'd14912:data <=32'hFFEEFFB3;
14'd14913:data <=32'hFFFBFFB4;14'd14914:data <=32'h000BFFA0;14'd14915:data <=32'h0026FF1F;
14'd14916:data <=32'h001FFEE9;14'd14917:data <=32'hFFE8FEE9;14'd14918:data <=32'hFFB3FEF8;
14'd14919:data <=32'hFF84FF14;14'd14920:data <=32'hFF61FF3A;14'd14921:data <=32'hFF48FF63;
14'd14922:data <=32'hFF3CFF8E;14'd14923:data <=32'hFF39FFB8;14'd14924:data <=32'hFF3EFFDF;
14'd14925:data <=32'hFF4C0003;14'd14926:data <=32'hFF610021;14'd14927:data <=32'hFF7D0037;
14'd14928:data <=32'hFF9B0044;14'd14929:data <=32'hFFBB0046;14'd14930:data <=32'hFFD6003C;
14'd14931:data <=32'hFFEA0029;14'd14932:data <=32'hFFF20013;14'd14933:data <=32'hFFF0FFFE;
14'd14934:data <=32'hFFE3FFEF;14'd14935:data <=32'hFFD2FFE8;14'd14936:data <=32'hFFC0FFEA;
14'd14937:data <=32'hFFB2FFF4;14'd14938:data <=32'hFFA90003;14'd14939:data <=32'hFFA70012;
14'd14940:data <=32'hFFA90022;14'd14941:data <=32'hFFAE002E;14'd14942:data <=32'hFFB70039;
14'd14943:data <=32'hFFC10041;14'd14944:data <=32'hFFCB0047;14'd14945:data <=32'hFFD6004B;
14'd14946:data <=32'hFFE3004B;14'd14947:data <=32'hFFEE0048;14'd14948:data <=32'hFFF70041;
14'd14949:data <=32'hFFFD0038;14'd14950:data <=32'hFFFD002E;14'd14951:data <=32'hFFF80026;
14'd14952:data <=32'hFFF00022;14'd14953:data <=32'hFFE60025;14'd14954:data <=32'hFFDD002C;
14'd14955:data <=32'hFFDA0038;14'd14956:data <=32'hFFDB0045;14'd14957:data <=32'hFFE30051;
14'd14958:data <=32'hFFED005A;14'd14959:data <=32'hFFF7005F;14'd14960:data <=32'h00010061;
14'd14961:data <=32'h00080062;14'd14962:data <=32'h000D0063;14'd14963:data <=32'h00120069;
14'd14964:data <=32'h001A0070;14'd14965:data <=32'h0024007A;14'd14966:data <=32'h00350082;
14'd14967:data <=32'h004A0088;14'd14968:data <=32'h00640088;14'd14969:data <=32'h007E0083;
14'd14970:data <=32'h00990079;14'd14971:data <=32'h00B40068;14'd14972:data <=32'h00CD0053;
14'd14973:data <=32'h00E60037;14'd14974:data <=32'h00FC0015;14'd14975:data <=32'h010DFFEA;
14'd14976:data <=32'h0058FFAD;14'd14977:data <=32'h0061FFAB;14'd14978:data <=32'h0079FFAD;
14'd14979:data <=32'h00F9FF9A;14'd14980:data <=32'h0106FF38;14'd14981:data <=32'h00D6FF08;
14'd14982:data <=32'h009AFEE7;14'd14983:data <=32'h005BFED8;14'd14984:data <=32'h001EFEDA;
14'd14985:data <=32'hFFE7FEE8;14'd14986:data <=32'hFFB9FEFF;14'd14987:data <=32'hFF92FF20;
14'd14988:data <=32'hFF74FF44;14'd14989:data <=32'hFF61FF6C;14'd14990:data <=32'hFF58FF96;
14'd14991:data <=32'hFF5AFFC0;14'd14992:data <=32'hFF66FFE4;14'd14993:data <=32'hFF7B0000;
14'd14994:data <=32'hFF950013;14'd14995:data <=32'hFFAF0019;14'd14996:data <=32'hFFC50016;
14'd14997:data <=32'hFFD4000E;14'd14998:data <=32'hFFDC0003;14'd14999:data <=32'hFFDCFFFA;
14'd15000:data <=32'hFFDAFFF5;14'd15001:data <=32'hFFD7FFF3;14'd15002:data <=32'hFFD5FFF4;
14'd15003:data <=32'hFFD6FFF5;14'd15004:data <=32'hFFD7FFF4;14'd15005:data <=32'hFFD7FFF2;
14'd15006:data <=32'hFFD5FFEE;14'd15007:data <=32'hFFD0FFEB;14'd15008:data <=32'hFFC8FFEA;
14'd15009:data <=32'hFFC0FFEC;14'd15010:data <=32'hFFB8FFF1;14'd15011:data <=32'hFFB1FFF8;
14'd15012:data <=32'hFFAC0002;14'd15013:data <=32'hFFA9000A;14'd15014:data <=32'hFFA70015;
14'd15015:data <=32'hFFA5001F;14'd15016:data <=32'hFFA5002A;14'd15017:data <=32'hFFA70038;
14'd15018:data <=32'hFFAB0047;14'd15019:data <=32'hFFB50055;14'd15020:data <=32'hFFC40060;
14'd15021:data <=32'hFFD60068;14'd15022:data <=32'hFFEA0068;14'd15023:data <=32'hFFFB0060;
14'd15024:data <=32'h00080052;14'd15025:data <=32'h000B0042;14'd15026:data <=32'h00060035;
14'd15027:data <=32'hFFFB002C;14'd15028:data <=32'hFFEA002D;14'd15029:data <=32'hFFDC0036;
14'd15030:data <=32'hFFD30047;14'd15031:data <=32'hFFCF005D;14'd15032:data <=32'hFFD30077;
14'd15033:data <=32'hFFE00090;14'd15034:data <=32'hFFF400A6;14'd15035:data <=32'h001000BA;
14'd15036:data <=32'h003300C7;14'd15037:data <=32'h005D00CF;14'd15038:data <=32'h008B00CB;
14'd15039:data <=32'h00BD00BB;14'd15040:data <=32'h008C0068;14'd15041:data <=32'h00B40062;
14'd15042:data <=32'h00C8005D;14'd15043:data <=32'h00CF0076;14'd15044:data <=32'h010A001F;
14'd15045:data <=32'h0106FFED;14'd15046:data <=32'h00F6FFC0;14'd15047:data <=32'h00DFFF9B;
14'd15048:data <=32'h00C3FF7E;14'd15049:data <=32'h00A6FF6B;14'd15050:data <=32'h008AFF5B;
14'd15051:data <=32'h006EFF51;14'd15052:data <=32'h0051FF4A;14'd15053:data <=32'h0034FF47;
14'd15054:data <=32'h0019FF49;14'd15055:data <=32'hFFFEFF52;14'd15056:data <=32'hFFE8FF5F;
14'd15057:data <=32'hFFD7FF6E;14'd15058:data <=32'hFFCBFF7C;14'd15059:data <=32'hFFC2FF8A;
14'd15060:data <=32'hFFBBFF95;14'd15061:data <=32'hFFB2FFA0;14'd15062:data <=32'hFFA9FFAC;
14'd15063:data <=32'hFFA1FFBC;14'd15064:data <=32'hFF9BFFCF;14'd15065:data <=32'hFF9BFFE6;
14'd15066:data <=32'hFFA3FFFC;14'd15067:data <=32'hFFB2000E;14'd15068:data <=32'hFFC7001A;
14'd15069:data <=32'hFFDE001D;14'd15070:data <=32'hFFF30016;14'd15071:data <=32'h00030009;
14'd15072:data <=32'h000DFFF6;14'd15073:data <=32'h000FFFE2;14'd15074:data <=32'h0009FFD0;
14'd15075:data <=32'hFFFEFFC0;14'd15076:data <=32'hFFEFFFB5;14'd15077:data <=32'hFFDDFFAD;
14'd15078:data <=32'hFFC6FFAA;14'd15079:data <=32'hFFB0FFAD;14'd15080:data <=32'hFF99FFB7;
14'd15081:data <=32'hFF85FFC6;14'd15082:data <=32'hFF75FFDD;14'd15083:data <=32'hFF6BFFF8;
14'd15084:data <=32'hFF6C0016;14'd15085:data <=32'hFF740032;14'd15086:data <=32'hFF850048;
14'd15087:data <=32'hFF9B0056;14'd15088:data <=32'hFFB0005A;14'd15089:data <=32'hFFC10058;
14'd15090:data <=32'hFFCD0051;14'd15091:data <=32'hFFD10049;14'd15092:data <=32'hFFCF0043;
14'd15093:data <=32'hFFCA0045;14'd15094:data <=32'hFFC4004A;14'd15095:data <=32'hFFC10055;
14'd15096:data <=32'hFFC10063;14'd15097:data <=32'hFFC50072;14'd15098:data <=32'hFFCE0082;
14'd15099:data <=32'hFFDA0090;14'd15100:data <=32'hFFEA009E;14'd15101:data <=32'hFFFE00AC;
14'd15102:data <=32'h001900B7;14'd15103:data <=32'h003800BC;14'd15104:data <=32'hFFD200D1;
14'd15105:data <=32'h000500FC;14'd15106:data <=32'h003A0101;14'd15107:data <=32'h0056008F;
14'd15108:data <=32'h008E0053;14'd15109:data <=32'h008D003B;14'd15110:data <=32'h00860028;
14'd15111:data <=32'h007C001B;14'd15112:data <=32'h00740016;14'd15113:data <=32'h00710016;
14'd15114:data <=32'h00740016;14'd15115:data <=32'h007C0012;14'd15116:data <=32'h0086000A;
14'd15117:data <=32'h0090FFFC;14'd15118:data <=32'h0096FFE9;14'd15119:data <=32'h0097FFD3;
14'd15120:data <=32'h0095FFBE;14'd15121:data <=32'h008FFFA8;14'd15122:data <=32'h0084FF91;
14'd15123:data <=32'h0075FF7C;14'd15124:data <=32'h0060FF67;14'd15125:data <=32'h0044FF55;
14'd15126:data <=32'h0022FF4B;14'd15127:data <=32'hFFFCFF49;14'd15128:data <=32'hFFD6FF54;
14'd15129:data <=32'hFFB4FF6C;14'd15130:data <=32'hFF9DFF8B;14'd15131:data <=32'hFF92FFAF;
14'd15132:data <=32'hFF94FFD3;14'd15133:data <=32'hFFA1FFF2;14'd15134:data <=32'hFFB40008;
14'd15135:data <=32'hFFCD0016;14'd15136:data <=32'hFFE60019;14'd15137:data <=32'hFFFB0015;
14'd15138:data <=32'h000E000C;14'd15139:data <=32'h001BFFFE;14'd15140:data <=32'h0024FFED;
14'd15141:data <=32'h0028FFD9;14'd15142:data <=32'h0027FFC5;14'd15143:data <=32'h001FFFB1;
14'd15144:data <=32'h0011FF9E;14'd15145:data <=32'hFFFDFF90;14'd15146:data <=32'hFFE6FF88;
14'd15147:data <=32'hFFCCFF88;14'd15148:data <=32'hFFB4FF8E;14'd15149:data <=32'hFFA0FF9A;
14'd15150:data <=32'hFF90FFA8;14'd15151:data <=32'hFF85FFB6;14'd15152:data <=32'hFF7CFFC4;
14'd15153:data <=32'hFF74FFD1;14'd15154:data <=32'hFF6BFFDC;14'd15155:data <=32'hFF5FFFEA;
14'd15156:data <=32'hFF53FFFD;14'd15157:data <=32'hFF490016;14'd15158:data <=32'hFF440035;
14'd15159:data <=32'hFF460057;14'd15160:data <=32'hFF520078;14'd15161:data <=32'hFF660098;
14'd15162:data <=32'hFF8100AF;14'd15163:data <=32'hFFA000C2;14'd15164:data <=32'hFFC100CE;
14'd15165:data <=32'hFFE200D2;14'd15166:data <=32'h000400D0;14'd15167:data <=32'h002400CA;
14'd15168:data <=32'hFF61005F;14'd15169:data <=32'hFF6800A0;14'd15170:data <=32'hFF9500D4;
14'd15171:data <=32'h004700AF;14'd15172:data <=32'h00820069;14'd15173:data <=32'h007C0045;
14'd15174:data <=32'h006D002A;14'd15175:data <=32'h00570017;14'd15176:data <=32'h00400013;
14'd15177:data <=32'h002D001A;14'd15178:data <=32'h00220029;14'd15179:data <=32'h00230039;
14'd15180:data <=32'h002C0047;14'd15181:data <=32'h003A004F;14'd15182:data <=32'h004D0052;
14'd15183:data <=32'h0061004F;14'd15184:data <=32'h00750046;14'd15185:data <=32'h00870038;
14'd15186:data <=32'h00970025;14'd15187:data <=32'h00A3000D;14'd15188:data <=32'h00AAFFEF;
14'd15189:data <=32'h00A9FFCE;14'd15190:data <=32'h009DFFAD;14'd15191:data <=32'h0086FF8F;
14'd15192:data <=32'h0069FF7A;14'd15193:data <=32'h0046FF70;14'd15194:data <=32'h0025FF71;
14'd15195:data <=32'h0007FF7C;14'd15196:data <=32'hFFF1FF8D;14'd15197:data <=32'hFFE4FF9F;
14'd15198:data <=32'hFFDEFFB3;14'd15199:data <=32'hFFDCFFC4;14'd15200:data <=32'hFFDEFFD1;
14'd15201:data <=32'hFFE1FFDC;14'd15202:data <=32'hFFE5FFE5;14'd15203:data <=32'hFFEBFFEF;
14'd15204:data <=32'hFFF3FFF7;14'd15205:data <=32'hFFFEFFFC;14'd15206:data <=32'h000BFFFE;
14'd15207:data <=32'h0019FFFB;14'd15208:data <=32'h0026FFF4;14'd15209:data <=32'h0031FFE7;
14'd15210:data <=32'h0038FFD7;14'd15211:data <=32'h003BFFC7;14'd15212:data <=32'h0039FFB4;
14'd15213:data <=32'h0035FFA2;14'd15214:data <=32'h002EFF8F;14'd15215:data <=32'h0022FF7B;
14'd15216:data <=32'h0011FF67;14'd15217:data <=32'hFFF9FF52;14'd15218:data <=32'hFFD9FF42;
14'd15219:data <=32'hFFAFFF38;14'd15220:data <=32'hFF81FF39;14'd15221:data <=32'hFF4FFF48;
14'd15222:data <=32'hFF21FF67;14'd15223:data <=32'hFEFCFF94;14'd15224:data <=32'hFEE3FFCA;
14'd15225:data <=32'hFED90004;14'd15226:data <=32'hFEDF003F;14'd15227:data <=32'hFEF30075;
14'd15228:data <=32'hFF1100A4;14'd15229:data <=32'hFF3700CA;14'd15230:data <=32'hFF6400E5;
14'd15231:data <=32'hFF9500F7;14'd15232:data <=32'hFF780037;14'd15233:data <=32'hFF6B005D;
14'd15234:data <=32'hFF6C0096;14'd15235:data <=32'hFFB500F9;14'd15236:data <=32'h000F00C8;
14'd15237:data <=32'h002700AE;14'd15238:data <=32'h00350092;14'd15239:data <=32'h00390079;
14'd15240:data <=32'h00350067;14'd15241:data <=32'h002F005E;14'd15242:data <=32'h002B005B;
14'd15243:data <=32'h002C005D;14'd15244:data <=32'h0032005D;14'd15245:data <=32'h003A005C;
14'd15246:data <=32'h00430058;14'd15247:data <=32'h004C0051;14'd15248:data <=32'h00530049;
14'd15249:data <=32'h00590041;14'd15250:data <=32'h005F0039;14'd15251:data <=32'h00640030;
14'd15252:data <=32'h006A0025;14'd15253:data <=32'h006E0017;14'd15254:data <=32'h006E0008;
14'd15255:data <=32'h006AFFF7;14'd15256:data <=32'h0061FFEA;14'd15257:data <=32'h0056FFE0;
14'd15258:data <=32'h004AFFDD;14'd15259:data <=32'h0040FFDD;14'd15260:data <=32'h003AFFE1;
14'd15261:data <=32'h0038FFE4;14'd15262:data <=32'h003BFFE4;14'd15263:data <=32'h003EFFE0;
14'd15264:data <=32'h003EFFD9;14'd15265:data <=32'h003BFFCF;14'd15266:data <=32'h0031FFC6;
14'd15267:data <=32'h0026FFC2;14'd15268:data <=32'h0019FFC1;14'd15269:data <=32'h000CFFC7;
14'd15270:data <=32'h0004FFD1;14'd15271:data <=32'h0001FFDD;14'd15272:data <=32'h0003FFE9;
14'd15273:data <=32'h0009FFF3;14'd15274:data <=32'h0013FFFA;14'd15275:data <=32'h0021FFFE;
14'd15276:data <=32'h0030FFFE;14'd15277:data <=32'h0041FFF9;14'd15278:data <=32'h0052FFEE;
14'd15279:data <=32'h0062FFDB;14'd15280:data <=32'h0071FFC2;14'd15281:data <=32'h0076FFA0;
14'd15282:data <=32'h0071FF79;14'd15283:data <=32'h005FFF50;14'd15284:data <=32'h003FFF2B;
14'd15285:data <=32'h0012FF11;14'd15286:data <=32'hFFDDFF05;14'd15287:data <=32'hFFA5FF07;
14'd15288:data <=32'hFF70FF19;14'd15289:data <=32'hFF43FF37;14'd15290:data <=32'hFF20FF5E;
14'd15291:data <=32'hFF08FF8B;14'd15292:data <=32'hFEFAFFB9;14'd15293:data <=32'hFEF4FFE7;
14'd15294:data <=32'hFEF80015;14'd15295:data <=32'hFF040040;14'd15296:data <=32'hFF240022;
14'd15297:data <=32'hFF1D004B;14'd15298:data <=32'hFF170068;14'd15299:data <=32'hFF030056;
14'd15300:data <=32'hFF470050;14'd15301:data <=32'hFF550061;14'd15302:data <=32'hFF620071;
14'd15303:data <=32'hFF6F0080;14'd15304:data <=32'hFF7A0091;14'd15305:data <=32'hFF8A00A5;
14'd15306:data <=32'hFF9F00B9;14'd15307:data <=32'hFFBC00CA;14'd15308:data <=32'hFFE000D5;
14'd15309:data <=32'h000700D7;14'd15310:data <=32'h002F00CB;14'd15311:data <=32'h005000B7;
14'd15312:data <=32'h006A009C;14'd15313:data <=32'h007A007D;14'd15314:data <=32'h0083005F;
14'd15315:data <=32'h00840041;14'd15316:data <=32'h007F0026;14'd15317:data <=32'h0075000E;
14'd15318:data <=32'h0067FFFA;14'd15319:data <=32'h0056FFEB;14'd15320:data <=32'h0040FFE2;
14'd15321:data <=32'h0028FFE1;14'd15322:data <=32'h0013FFE9;14'd15323:data <=32'h0004FFF7;
14'd15324:data <=32'hFFFE000B;14'd15325:data <=32'h00000020;14'd15326:data <=32'h000D0030;
14'd15327:data <=32'h001E0039;14'd15328:data <=32'h0032003A;14'd15329:data <=32'h00440033;
14'd15330:data <=32'h00510026;14'd15331:data <=32'h00560016;14'd15332:data <=32'h00560007;
14'd15333:data <=32'h0053FFFB;14'd15334:data <=32'h004EFFF3;14'd15335:data <=32'h0047FFEE;
14'd15336:data <=32'h0042FFEB;14'd15337:data <=32'h003EFFEA;14'd15338:data <=32'h003CFFEA;
14'd15339:data <=32'h003BFFEA;14'd15340:data <=32'h003BFFEB;14'd15341:data <=32'h003EFFEE;
14'd15342:data <=32'h0044FFED;14'd15343:data <=32'h004DFFEC;14'd15344:data <=32'h0059FFE5;
14'd15345:data <=32'h0064FFD8;14'd15346:data <=32'h006DFFC5;14'd15347:data <=32'h006FFFAC;
14'd15348:data <=32'h0069FF90;14'd15349:data <=32'h005BFF75;14'd15350:data <=32'h0044FF61;
14'd15351:data <=32'h0028FF53;14'd15352:data <=32'h000BFF4E;14'd15353:data <=32'hFFF1FF50;
14'd15354:data <=32'hFFD9FF56;14'd15355:data <=32'hFFC8FF5D;14'd15356:data <=32'hFFB7FF65;
14'd15357:data <=32'hFFA8FF6C;14'd15358:data <=32'hFF97FF73;14'd15359:data <=32'hFF85FF7C;
14'd15360:data <=32'hFF1DFF66;14'd15361:data <=32'hFEF7FF8C;14'd15362:data <=32'hFEF3FFB1;
14'd15363:data <=32'hFF60FF83;14'd15364:data <=32'hFF7CFF6D;14'd15365:data <=32'hFF60FF77;
14'd15366:data <=32'hFF41FF88;14'd15367:data <=32'hFF23FFA1;14'd15368:data <=32'hFF07FFC6;
14'd15369:data <=32'hFEF3FFF3;14'd15370:data <=32'hFEEB0029;14'd15371:data <=32'hFEF40064;
14'd15372:data <=32'hFF0D009A;14'd15373:data <=32'hFF3400C9;14'd15374:data <=32'hFF6800E8;
14'd15375:data <=32'hFFA000F9;14'd15376:data <=32'hFFD600FA;14'd15377:data <=32'h000800EE;
14'd15378:data <=32'h003300D8;14'd15379:data <=32'h005400BB;14'd15380:data <=32'h006D009A;
14'd15381:data <=32'h007C0075;14'd15382:data <=32'h0083004F;14'd15383:data <=32'h007F002B;
14'd15384:data <=32'h0071000A;14'd15385:data <=32'h005AFFF0;14'd15386:data <=32'h0040FFE1;
14'd15387:data <=32'h0022FFDC;14'd15388:data <=32'h0007FFE2;14'd15389:data <=32'hFFF4FFF0;
14'd15390:data <=32'hFFE80004;14'd15391:data <=32'hFFE50017;14'd15392:data <=32'hFFE90028;
14'd15393:data <=32'hFFF00034;14'd15394:data <=32'hFFF9003C;14'd15395:data <=32'h00010042;
14'd15396:data <=32'h00090047;14'd15397:data <=32'h0011004C;14'd15398:data <=32'h001A0052;
14'd15399:data <=32'h00270056;14'd15400:data <=32'h0036005A;14'd15401:data <=32'h00480059;
14'd15402:data <=32'h005A0054;14'd15403:data <=32'h006C0049;14'd15404:data <=32'h007C003A;
14'd15405:data <=32'h0087002A;14'd15406:data <=32'h00900017;14'd15407:data <=32'h00950003;
14'd15408:data <=32'h0098FFEF;14'd15409:data <=32'h0098FFD8;14'd15410:data <=32'h0094FFC0;
14'd15411:data <=32'h008BFFA8;14'd15412:data <=32'h007BFF92;14'd15413:data <=32'h0065FF80;
14'd15414:data <=32'h004AFF75;14'd15415:data <=32'h002EFF73;14'd15416:data <=32'h0015FF7B;
14'd15417:data <=32'h0002FF88;14'd15418:data <=32'hFFFAFF9A;14'd15419:data <=32'hFFFAFFA9;
14'd15420:data <=32'h0002FFB3;14'd15421:data <=32'h000DFFB4;14'd15422:data <=32'h0016FFAE;
14'd15423:data <=32'h001BFFA0;14'd15424:data <=32'hFFEEFF1F;14'd15425:data <=32'hFFC4FF16;
14'd15426:data <=32'hFFA5FF30;14'd15427:data <=32'hFFEFFF8B;14'd15428:data <=32'h0018FF5E;
14'd15429:data <=32'h0000FF4A;14'd15430:data <=32'hFFE0FF3A;14'd15431:data <=32'hFFBAFF32;
14'd15432:data <=32'hFF8DFF35;14'd15433:data <=32'hFF5EFF45;14'd15434:data <=32'hFF34FF64;
14'd15435:data <=32'hFF14FF91;14'd15436:data <=32'hFF02FFC4;14'd15437:data <=32'hFEFFFFF9;
14'd15438:data <=32'hFF0B002B;14'd15439:data <=32'hFF220055;14'd15440:data <=32'hFF3F0075;
14'd15441:data <=32'hFF5F008B;14'd15442:data <=32'hFF81009A;14'd15443:data <=32'hFFA200A3;
14'd15444:data <=32'hFFC100A4;14'd15445:data <=32'hFFE000A0;14'd15446:data <=32'hFFFD0098;
14'd15447:data <=32'h00150088;14'd15448:data <=32'h00270073;14'd15449:data <=32'h0033005D;
14'd15450:data <=32'h00370046;14'd15451:data <=32'h00340032;14'd15452:data <=32'h002D0022;
14'd15453:data <=32'h00250017;14'd15454:data <=32'h001C0010;14'd15455:data <=32'h0015000B;
14'd15456:data <=32'h000E0005;14'd15457:data <=32'h00050001;14'd15458:data <=32'hFFFAFFFD;
14'd15459:data <=32'hFFEBFFFC;14'd15460:data <=32'hFFDA0002;14'd15461:data <=32'hFFC9000E;
14'd15462:data <=32'hFFBC0022;14'd15463:data <=32'hFFB5003C;14'd15464:data <=32'hFFB8005A;
14'd15465:data <=32'hFFC40078;14'd15466:data <=32'hFFDA0091;14'd15467:data <=32'hFFF800A3;
14'd15468:data <=32'h001B00AE;14'd15469:data <=32'h003F00AF;14'd15470:data <=32'h006300A8;
14'd15471:data <=32'h00860098;14'd15472:data <=32'h00A40081;14'd15473:data <=32'h00BE0064;
14'd15474:data <=32'h00D10040;14'd15475:data <=32'h00DB0017;14'd15476:data <=32'h00DAFFEC;
14'd15477:data <=32'h00CCFFC3;14'd15478:data <=32'h00B5FF9F;14'd15479:data <=32'h0095FF87;
14'd15480:data <=32'h0071FF7B;14'd15481:data <=32'h0050FF7B;14'd15482:data <=32'h0035FF86;
14'd15483:data <=32'h0025FF95;14'd15484:data <=32'h001FFFA5;14'd15485:data <=32'h0020FFB1;
14'd15486:data <=32'h0025FFB7;14'd15487:data <=32'h002EFFB6;14'd15488:data <=32'h0050FFAE;
14'd15489:data <=32'h0054FF99;14'd15490:data <=32'h0040FF87;14'd15491:data <=32'h0004FF8D;
14'd15492:data <=32'h0030FF6E;14'd15493:data <=32'h0021FF64;14'd15494:data <=32'h000FFF5C;
14'd15495:data <=32'hFFFAFF55;14'd15496:data <=32'hFFE0FF52;14'd15497:data <=32'hFFC3FF55;
14'd15498:data <=32'hFFA5FF61;14'd15499:data <=32'hFF8DFF75;14'd15500:data <=32'hFF7BFF90;
14'd15501:data <=32'hFF73FFAB;14'd15502:data <=32'hFF74FFC6;14'd15503:data <=32'hFF7AFFDB;
14'd15504:data <=32'hFF83FFEB;14'd15505:data <=32'hFF8BFFF2;14'd15506:data <=32'hFF90FFF9;
14'd15507:data <=32'hFF91FFFF;14'd15508:data <=32'hFF910006;14'd15509:data <=32'hFF910011;
14'd15510:data <=32'hFF93001D;14'd15511:data <=32'hFF980029;14'd15512:data <=32'hFFA00034;
14'd15513:data <=32'hFFA9003D;14'd15514:data <=32'hFFB40045;14'd15515:data <=32'hFFBE004B;
14'd15516:data <=32'hFFCB0051;14'd15517:data <=32'hFFD80056;14'd15518:data <=32'hFFE80057;
14'd15519:data <=32'hFFFA0054;14'd15520:data <=32'h000B004A;14'd15521:data <=32'h0018003B;
14'd15522:data <=32'h001F0024;14'd15523:data <=32'h001E000D;14'd15524:data <=32'h0012FFF7;
14'd15525:data <=32'hFFFDFFE8;14'd15526:data <=32'hFFE3FFE2;14'd15527:data <=32'hFFC7FFE7;
14'd15528:data <=32'hFFADFFF6;14'd15529:data <=32'hFF9B000F;14'd15530:data <=32'hFF92002C;
14'd15531:data <=32'hFF91004C;14'd15532:data <=32'hFF9A006A;14'd15533:data <=32'hFFAA0086;
14'd15534:data <=32'hFFC0009E;14'd15535:data <=32'hFFDB00B1;14'd15536:data <=32'hFFFB00BD;
14'd15537:data <=32'h001D00C3;14'd15538:data <=32'h004200C2;14'd15539:data <=32'h006500B5;
14'd15540:data <=32'h008600A1;14'd15541:data <=32'h00A00085;14'd15542:data <=32'h00AE0066;
14'd15543:data <=32'h00B60048;14'd15544:data <=32'h00B5002D;14'd15545:data <=32'h00B10017;
14'd15546:data <=32'h00AB0006;14'd15547:data <=32'h00A8FFF9;14'd15548:data <=32'h00A8FFEC;
14'd15549:data <=32'h00ABFFDC;14'd15550:data <=32'h00ACFFC9;14'd15551:data <=32'h00AAFFB2;
14'd15552:data <=32'h0023FFDF;14'd15553:data <=32'h0035FFE7;14'd15554:data <=32'h004DFFDC;
14'd15555:data <=32'h0087FF6D;14'd15556:data <=32'h00A0FF3F;14'd15557:data <=32'h007AFF2A;
14'd15558:data <=32'h0051FF1E;14'd15559:data <=32'h0028FF1C;14'd15560:data <=32'hFFFFFF20;
14'd15561:data <=32'hFFD7FF2C;14'd15562:data <=32'hFFB4FF43;14'd15563:data <=32'hFF99FF63;
14'd15564:data <=32'hFF88FF88;14'd15565:data <=32'hFF85FFAE;14'd15566:data <=32'hFF8FFFD0;
14'd15567:data <=32'hFFA0FFE8;14'd15568:data <=32'hFFB9FFF5;14'd15569:data <=32'hFFD0FFF8;
14'd15570:data <=32'hFFE0FFF0;14'd15571:data <=32'hFFE8FFE4;14'd15572:data <=32'hFFEAFFD6;
14'd15573:data <=32'hFFE3FFCA;14'd15574:data <=32'hFFDAFFC4;14'd15575:data <=32'hFFCDFFC1;
14'd15576:data <=32'hFFC1FFC2;14'd15577:data <=32'hFFB3FFC6;14'd15578:data <=32'hFFA8FFCE;
14'd15579:data <=32'hFF9DFFDB;14'd15580:data <=32'hFF95FFEA;14'd15581:data <=32'hFF91FFFD;
14'd15582:data <=32'hFF930012;14'd15583:data <=32'hFF9C0025;14'd15584:data <=32'hFFAD0035;
14'd15585:data <=32'hFFBF003C;14'd15586:data <=32'hFFD4003C;14'd15587:data <=32'hFFE50034;
14'd15588:data <=32'hFFF00027;14'd15589:data <=32'hFFF30017;14'd15590:data <=32'hFFEE0009;
14'd15591:data <=32'hFFE40000;14'd15592:data <=32'hFFD8FFFD;14'd15593:data <=32'hFFCCFFFE;
14'd15594:data <=32'hFFC20005;14'd15595:data <=32'hFFBA000D;14'd15596:data <=32'hFFB50016;
14'd15597:data <=32'hFFB10020;14'd15598:data <=32'hFFAE002A;14'd15599:data <=32'hFFAA0035;
14'd15600:data <=32'hFFA90043;14'd15601:data <=32'hFFA90053;14'd15602:data <=32'hFFAE0064;
14'd15603:data <=32'hFFB70077;14'd15604:data <=32'hFFC20087;14'd15605:data <=32'hFFD20094;
14'd15606:data <=32'hFFE200A0;14'd15607:data <=32'hFFF300AA;14'd15608:data <=32'h000700B5;
14'd15609:data <=32'h001D00BE;14'd15610:data <=32'h003900C8;14'd15611:data <=32'h005B00CF;
14'd15612:data <=32'h008400CD;14'd15613:data <=32'h00B100C0;14'd15614:data <=32'h00DD00A7;
14'd15615:data <=32'h0104007F;14'd15616:data <=32'h005EFFF9;14'd15617:data <=32'h00660000;
14'd15618:data <=32'h007C0012;14'd15619:data <=32'h01070029;14'd15620:data <=32'h013BFFDC;
14'd15621:data <=32'h0129FFA2;14'd15622:data <=32'h010BFF6E;14'd15623:data <=32'h00E3FF46;
14'd15624:data <=32'h00B4FF26;14'd15625:data <=32'h007EFF12;14'd15626:data <=32'h0047FF0D;
14'd15627:data <=32'h0012FF16;14'd15628:data <=32'hFFE5FF2D;14'd15629:data <=32'hFFC3FF4F;
14'd15630:data <=32'hFFAFFF75;14'd15631:data <=32'hFFAAFF9A;14'd15632:data <=32'hFFB0FFB8;
14'd15633:data <=32'hFFBEFFCE;14'd15634:data <=32'hFFCDFFDA;14'd15635:data <=32'hFFDBFFDF;
14'd15636:data <=32'hFFE6FFDE;14'd15637:data <=32'hFFECFFDB;14'd15638:data <=32'hFFEEFFD8;
14'd15639:data <=32'hFFF0FFD6;14'd15640:data <=32'hFFF0FFD3;14'd15641:data <=32'hFFF1FFCE;
14'd15642:data <=32'hFFEEFFCA;14'd15643:data <=32'hFFEAFFC5;14'd15644:data <=32'hFFE2FFC2;
14'd15645:data <=32'hFFD9FFC2;14'd15646:data <=32'hFFD0FFC5;14'd15647:data <=32'hFFC8FFCB;
14'd15648:data <=32'hFFC4FFD2;14'd15649:data <=32'hFFC3FFD9;14'd15650:data <=32'hFFC3FFDD;
14'd15651:data <=32'hFFC4FFE0;14'd15652:data <=32'hFFC2FFDF;14'd15653:data <=32'hFFBDFFE0;
14'd15654:data <=32'hFFB5FFE1;14'd15655:data <=32'hFFADFFE8;14'd15656:data <=32'hFFA5FFF4;
14'd15657:data <=32'hFFA10001;14'd15658:data <=32'hFFA30010;14'd15659:data <=32'hFFAB001E;
14'd15660:data <=32'hFFB60027;14'd15661:data <=32'hFFC30029;14'd15662:data <=32'hFFCE0026;
14'd15663:data <=32'hFFD4001F;14'd15664:data <=32'hFFD50016;14'd15665:data <=32'hFFD0000E;
14'd15666:data <=32'hFFC80009;14'd15667:data <=32'hFFBC0008;14'd15668:data <=32'hFFAE000B;
14'd15669:data <=32'hFF9E0013;14'd15670:data <=32'hFF8F0020;14'd15671:data <=32'hFF810034;
14'd15672:data <=32'hFF75004F;14'd15673:data <=32'hFF700071;14'd15674:data <=32'hFF75009A;
14'd15675:data <=32'hFF8500C5;14'd15676:data <=32'hFFA600F0;14'd15677:data <=32'hFFD50110;
14'd15678:data <=32'h000F0125;14'd15679:data <=32'h00500127;14'd15680:data <=32'h004100A0;
14'd15681:data <=32'h006100AC;14'd15682:data <=32'h007000B6;14'd15683:data <=32'h007300E7;
14'd15684:data <=32'h00CF00B4;14'd15685:data <=32'h00E6008B;14'd15686:data <=32'h00F50060;
14'd15687:data <=32'h00FB0035;14'd15688:data <=32'h00F80009;14'd15689:data <=32'h00EEFFE0;
14'd15690:data <=32'h00DAFFBB;14'd15691:data <=32'h00BFFF9E;14'd15692:data <=32'h00A0FF8A;
14'd15693:data <=32'h0082FF80;14'd15694:data <=32'h0068FF7E;14'd15695:data <=32'h0053FF81;
14'd15696:data <=32'h0042FF83;14'd15697:data <=32'h0037FF85;14'd15698:data <=32'h002AFF83;
14'd15699:data <=32'h001CFF82;14'd15700:data <=32'h000AFF82;14'd15701:data <=32'hFFF7FF86;
14'd15702:data <=32'hFFE5FF90;14'd15703:data <=32'hFFD7FFA0;14'd15704:data <=32'hFFCEFFB3;
14'd15705:data <=32'hFFCBFFC6;14'd15706:data <=32'hFFCFFFD8;14'd15707:data <=32'hFFD6FFE5;
14'd15708:data <=32'hFFE2FFEE;14'd15709:data <=32'hFFEDFFF2;14'd15710:data <=32'hFFF8FFF5;
14'd15711:data <=32'h0004FFF2;14'd15712:data <=32'h000EFFEC;14'd15713:data <=32'h0017FFE3;
14'd15714:data <=32'h001EFFD6;14'd15715:data <=32'h0020FFC4;14'd15716:data <=32'h001BFFB0;
14'd15717:data <=32'h000EFF9E;14'd15718:data <=32'hFFFAFF90;14'd15719:data <=32'hFFE0FF8A;
14'd15720:data <=32'hFFC3FF8B;14'd15721:data <=32'hFFABFF97;14'd15722:data <=32'hFF97FFAB;
14'd15723:data <=32'hFF8BFFC3;14'd15724:data <=32'hFF89FFDB;14'd15725:data <=32'hFF8FFFEF;
14'd15726:data <=32'hFF98FFFD;14'd15727:data <=32'hFFA40005;14'd15728:data <=32'hFFAD0008;
14'd15729:data <=32'hFFB40008;14'd15730:data <=32'hFFB70006;14'd15731:data <=32'hFFB70002;
14'd15732:data <=32'hFFB4FFFF;14'd15733:data <=32'hFFAEFFFD;14'd15734:data <=32'hFFA4FFFD;
14'd15735:data <=32'hFF96FFFF;14'd15736:data <=32'hFF860007;14'd15737:data <=32'hFF760017;
14'd15738:data <=32'hFF66002F;14'd15739:data <=32'hFF5F004F;14'd15740:data <=32'hFF610075;
14'd15741:data <=32'hFF6F009C;14'd15742:data <=32'hFF8900BE;14'd15743:data <=32'hFFAE00D7;
14'd15744:data <=32'hFF6900B3;14'd15745:data <=32'hFF8300EB;14'd15746:data <=32'hFFA70101;
14'd15747:data <=32'hFFD500B1;14'd15748:data <=32'h0020009C;14'd15749:data <=32'h002D0094;
14'd15750:data <=32'h0037008D;14'd15751:data <=32'h00400087;14'd15752:data <=32'h004D0083;
14'd15753:data <=32'h0059007B;14'd15754:data <=32'h00660074;14'd15755:data <=32'h00710069;
14'd15756:data <=32'h007C005F;14'd15757:data <=32'h00870055;14'd15758:data <=32'h00940049;
14'd15759:data <=32'h00A2003B;14'd15760:data <=32'h00B10027;14'd15761:data <=32'h00BD000B;
14'd15762:data <=32'h00C3FFEA;14'd15763:data <=32'h00BFFFC5;14'd15764:data <=32'h00AFFF9E;
14'd15765:data <=32'h0094FF7F;14'd15766:data <=32'h0070FF68;14'd15767:data <=32'h0049FF5E;
14'd15768:data <=32'h0022FF61;14'd15769:data <=32'h0001FF6E;14'd15770:data <=32'hFFE6FF82;
14'd15771:data <=32'hFFD4FF9A;14'd15772:data <=32'hFFC9FFB4;14'd15773:data <=32'hFFC7FFCE;
14'd15774:data <=32'hFFCBFFE6;14'd15775:data <=32'hFFD5FFFC;14'd15776:data <=32'hFFE6000D;
14'd15777:data <=32'hFFFB0017;14'd15778:data <=32'h0013001A;14'd15779:data <=32'h002C0013;
14'd15780:data <=32'h00410004;14'd15781:data <=32'h004FFFEE;14'd15782:data <=32'h0055FFD2;
14'd15783:data <=32'h0050FFB8;14'd15784:data <=32'h0043FFA1;14'd15785:data <=32'h0031FF90;
14'd15786:data <=32'h001CFF86;14'd15787:data <=32'h0009FF82;14'd15788:data <=32'hFFF7FF82;
14'd15789:data <=32'hFFE9FF84;14'd15790:data <=32'hFFDCFF85;14'd15791:data <=32'hFFD0FF85;
14'd15792:data <=32'hFFC1FF85;14'd15793:data <=32'hFFB0FF87;14'd15794:data <=32'hFF9DFF8C;
14'd15795:data <=32'hFF8AFF95;14'd15796:data <=32'hFF78FFA4;14'd15797:data <=32'hFF68FFB5;
14'd15798:data <=32'hFF5CFFC9;14'd15799:data <=32'hFF53FFDE;14'd15800:data <=32'hFF4CFFF4;
14'd15801:data <=32'hFF48000C;14'd15802:data <=32'hFF470027;14'd15803:data <=32'hFF4A0044;
14'd15804:data <=32'hFF550063;14'd15805:data <=32'hFF67007F;14'd15806:data <=32'hFF810096;
14'd15807:data <=32'hFFA100A5;14'd15808:data <=32'hFF260002;14'd15809:data <=32'hFF0F003C;
14'd15810:data <=32'hFF1E0079;14'd15811:data <=32'hFFC7008C;14'd15812:data <=32'h000D006D;
14'd15813:data <=32'h000D0058;14'd15814:data <=32'h0006004A;14'd15815:data <=32'hFFFB0043;
14'd15816:data <=32'hFFF10045;14'd15817:data <=32'hFFEA004B;14'd15818:data <=32'hFFE60055;
14'd15819:data <=32'hFFE50062;14'd15820:data <=32'hFFEA0071;14'd15821:data <=32'hFFF40083;
14'd15822:data <=32'h00050094;14'd15823:data <=32'h001E00A1;14'd15824:data <=32'h003F00A7;
14'd15825:data <=32'h006400A3;14'd15826:data <=32'h00890092;14'd15827:data <=32'h00A80075;
14'd15828:data <=32'h00BE004F;14'd15829:data <=32'h00C60023;14'd15830:data <=32'h00C1FFFA;
14'd15831:data <=32'h00B1FFD5;14'd15832:data <=32'h009AFFBA;14'd15833:data <=32'h007EFFA7;
14'd15834:data <=32'h0063FF9D;14'd15835:data <=32'h0048FF99;14'd15836:data <=32'h0030FF9B;
14'd15837:data <=32'h001BFFA0;14'd15838:data <=32'h0007FFAB;14'd15839:data <=32'hFFF7FFB9;
14'd15840:data <=32'hFFEDFFCB;14'd15841:data <=32'hFFE9FFDF;14'd15842:data <=32'hFFECFFF2;
14'd15843:data <=32'hFFF50003;14'd15844:data <=32'h0002000F;14'd15845:data <=32'h00130015;
14'd15846:data <=32'h00230016;14'd15847:data <=32'h00320011;14'd15848:data <=32'h003D000A;
14'd15849:data <=32'h00480002;14'd15850:data <=32'h0052FFF9;14'd15851:data <=32'h005BFFEF;
14'd15852:data <=32'h0066FFE1;14'd15853:data <=32'h0070FFCF;14'd15854:data <=32'h0078FFB6;
14'd15855:data <=32'h0079FF97;14'd15856:data <=32'h0073FF74;14'd15857:data <=32'h0060FF51;
14'd15858:data <=32'h0043FF31;14'd15859:data <=32'h001BFF1B;14'd15860:data <=32'hFFEEFF0E;
14'd15861:data <=32'hFFBEFF0D;14'd15862:data <=32'hFF8FFF17;14'd15863:data <=32'hFF62FF2C;
14'd15864:data <=32'hFF3BFF49;14'd15865:data <=32'hFF1AFF6E;14'd15866:data <=32'hFF01FF9A;
14'd15867:data <=32'hFEF2FFCD;14'd15868:data <=32'hFEEF0002;14'd15869:data <=32'hFEFB0037;
14'd15870:data <=32'hFF150068;14'd15871:data <=32'hFF3B008D;14'd15872:data <=32'hFF70FFCB;
14'd15873:data <=32'hFF51FFE2;14'd15874:data <=32'hFF36000F;14'd15875:data <=32'hFF59008A;
14'd15876:data <=32'hFFB1007D;14'd15877:data <=32'hFFC40071;14'd15878:data <=32'hFFCF0066;
14'd15879:data <=32'hFFD3005C;14'd15880:data <=32'hFFD50057;14'd15881:data <=32'hFFD60054;
14'd15882:data <=32'hFFD70054;14'd15883:data <=32'hFFD80056;14'd15884:data <=32'hFFD7005A;
14'd15885:data <=32'hFFD80060;14'd15886:data <=32'hFFDC006A;14'd15887:data <=32'hFFE40076;
14'd15888:data <=32'hFFF20082;14'd15889:data <=32'h0006008A;14'd15890:data <=32'h001E008C;
14'd15891:data <=32'h00370085;14'd15892:data <=32'h004D0076;14'd15893:data <=32'h005C0063;
14'd15894:data <=32'h0063004E;14'd15895:data <=32'h0063003A;14'd15896:data <=32'h0060002B;
14'd15897:data <=32'h005B0020;14'd15898:data <=32'h0057001A;14'd15899:data <=32'h00540013;
14'd15900:data <=32'h0054000D;14'd15901:data <=32'h00530005;14'd15902:data <=32'h0050FFFC;
14'd15903:data <=32'h004CFFF2;14'd15904:data <=32'h0044FFEA;14'd15905:data <=32'h003BFFE5;
14'd15906:data <=32'h0031FFE3;14'd15907:data <=32'h0029FFE4;14'd15908:data <=32'h0021FFE6;
14'd15909:data <=32'h001AFFEA;14'd15910:data <=32'h0014FFF0;14'd15911:data <=32'h000FFFF6;
14'd15912:data <=32'h000B0001;14'd15913:data <=32'h000C000D;14'd15914:data <=32'h0010001C;
14'd15915:data <=32'h001C002C;14'd15916:data <=32'h002F0038;14'd15917:data <=32'h004C003F;
14'd15918:data <=32'h006D003B;14'd15919:data <=32'h008E0029;14'd15920:data <=32'h00AB000D;
14'd15921:data <=32'h00C0FFE5;14'd15922:data <=32'h00C7FFB6;14'd15923:data <=32'h00C1FF85;
14'd15924:data <=32'h00ADFF56;14'd15925:data <=32'h008EFF2F;14'd15926:data <=32'h0066FF0F;
14'd15927:data <=32'h0038FEF9;14'd15928:data <=32'h0007FEEF;14'd15929:data <=32'hFFD3FEED;
14'd15930:data <=32'hFFA0FEF7;14'd15931:data <=32'hFF70FF0E;14'd15932:data <=32'hFF46FF30;
14'd15933:data <=32'hFF25FF5A;14'd15934:data <=32'hFF12FF8B;14'd15935:data <=32'hFF0DFFBD;
14'd15936:data <=32'hFF51FFB3;14'd15937:data <=32'hFF40FFCA;14'd15938:data <=32'hFF2CFFD6;
14'd15939:data <=32'hFF0FFFC1;14'd15940:data <=32'hFF49FFD0;14'd15941:data <=32'hFF45FFE2;
14'd15942:data <=32'hFF3FFFF6;14'd15943:data <=32'hFF3B000E;14'd15944:data <=32'hFF3C002A;
14'd15945:data <=32'hFF440048;14'd15946:data <=32'hFF530065;14'd15947:data <=32'hFF68007B;
14'd15948:data <=32'hFF81008C;14'd15949:data <=32'hFF9B0099;14'd15950:data <=32'hFFB500A0;
14'd15951:data <=32'hFFCF00A3;14'd15952:data <=32'hFFEB00A3;14'd15953:data <=32'h0005009C;
14'd15954:data <=32'h001F0090;14'd15955:data <=32'h0035007D;14'd15956:data <=32'h00440064;
14'd15957:data <=32'h004A0049;14'd15958:data <=32'h0045002F;14'd15959:data <=32'h0038001A;
14'd15960:data <=32'h0026000E;14'd15961:data <=32'h0012000C;14'd15962:data <=32'h00030013;
14'd15963:data <=32'hFFFA0020;14'd15964:data <=32'hFFF8002D;14'd15965:data <=32'hFFFD003A;
14'd15966:data <=32'h00070042;14'd15967:data <=32'h00120046;14'd15968:data <=32'h001E0047;
14'd15969:data <=32'h00290044;14'd15970:data <=32'h0032003E;14'd15971:data <=32'h003A0037;
14'd15972:data <=32'h003F002E;14'd15973:data <=32'h00430024;14'd15974:data <=32'h0042001A;
14'd15975:data <=32'h003F0010;14'd15976:data <=32'h00380009;14'd15977:data <=32'h002E0007;
14'd15978:data <=32'h0024000B;14'd15979:data <=32'h001D0014;14'd15980:data <=32'h001C0022;
14'd15981:data <=32'h00240032;14'd15982:data <=32'h0034003E;14'd15983:data <=32'h004B0043;
14'd15984:data <=32'h00660041;14'd15985:data <=32'h007E0033;14'd15986:data <=32'h0093001E;
14'd15987:data <=32'h00A00004;14'd15988:data <=32'h00A6FFE7;14'd15989:data <=32'h00A5FFCA;
14'd15990:data <=32'h00A0FFAF;14'd15991:data <=32'h0096FF97;14'd15992:data <=32'h0089FF7F;
14'd15993:data <=32'h0078FF6A;14'd15994:data <=32'h0063FF57;14'd15995:data <=32'h004BFF47;
14'd15996:data <=32'h002FFF3C;14'd15997:data <=32'h0013FF38;14'd15998:data <=32'hFFF7FF39;
14'd15999:data <=32'hFFDFFF3F;14'd16000:data <=32'hFF8AFF22;14'd16001:data <=32'hFF66FF34;
14'd16002:data <=32'hFF5EFF48;14'd16003:data <=32'hFFCDFF2C;14'd16004:data <=32'hFFE9FF1C;
14'd16005:data <=32'hFFC0FF13;14'd16006:data <=32'hFF91FF14;14'd16007:data <=32'hFF5FFF23;
14'd16008:data <=32'hFF31FF41;14'd16009:data <=32'hFF0AFF6C;14'd16010:data <=32'hFEF2FFA0;
14'd16011:data <=32'hFEE9FFD7;14'd16012:data <=32'hFEEC000D;14'd16013:data <=32'hFEFB003F;
14'd16014:data <=32'hFF14006B;14'd16015:data <=32'hFF350091;14'd16016:data <=32'hFF5D00AE;
14'd16017:data <=32'hFF8A00C0;14'd16018:data <=32'hFFB900C7;14'd16019:data <=32'hFFE900C1;
14'd16020:data <=32'h001300AD;14'd16021:data <=32'h0032008F;14'd16022:data <=32'h0047006A;
14'd16023:data <=32'h004B0044;14'd16024:data <=32'h00440023;14'd16025:data <=32'h0033000B;
14'd16026:data <=32'h001EFFFD;14'd16027:data <=32'h0008FFF8;14'd16028:data <=32'hFFF6FFFA;
14'd16029:data <=32'hFFE90002;14'd16030:data <=32'hFFE0000B;14'd16031:data <=32'hFFDA0015;
14'd16032:data <=32'hFFD60020;14'd16033:data <=32'hFFD4002A;14'd16034:data <=32'hFFD50036;
14'd16035:data <=32'hFFD80042;14'd16036:data <=32'hFFDF004D;14'd16037:data <=32'hFFE80057;
14'd16038:data <=32'hFFF5005D;14'd16039:data <=32'h00010062;14'd16040:data <=32'h000D0063;
14'd16041:data <=32'h00180062;14'd16042:data <=32'h00210061;14'd16043:data <=32'h002A0061;
14'd16044:data <=32'h00340062;14'd16045:data <=32'h00400062;14'd16046:data <=32'h00510061;
14'd16047:data <=32'h0063005A;14'd16048:data <=32'h0075004E;14'd16049:data <=32'h0084003C;
14'd16050:data <=32'h008D0025;14'd16051:data <=32'h008F000C;14'd16052:data <=32'h0089FFF6;
14'd16053:data <=32'h007EFFE4;14'd16054:data <=32'h0070FFDA;14'd16055:data <=32'h0063FFD5;
14'd16056:data <=32'h005AFFD5;14'd16057:data <=32'h0056FFD7;14'd16058:data <=32'h0056FFD8;
14'd16059:data <=32'h0058FFD8;14'd16060:data <=32'h005CFFD5;14'd16061:data <=32'h0062FFCF;
14'd16062:data <=32'h0069FFC7;14'd16063:data <=32'h0070FFBB;14'd16064:data <=32'h005FFF39;
14'd16065:data <=32'h0046FF25;14'd16066:data <=32'h002DFF2F;14'd16067:data <=32'h0068FF94;
14'd16068:data <=32'h00A0FF6C;14'd16069:data <=32'h008BFF40;14'd16070:data <=32'h0069FF18;
14'd16071:data <=32'h003BFEFB;14'd16072:data <=32'h0003FEED;14'd16073:data <=32'hFFCAFEEF;
14'd16074:data <=32'hFF95FF00;14'd16075:data <=32'hFF68FF1D;14'd16076:data <=32'hFF44FF42;
14'd16077:data <=32'hFF2AFF6C;14'd16078:data <=32'hFF1AFF98;14'd16079:data <=32'hFF12FFC5;
14'd16080:data <=32'hFF15FFF3;14'd16081:data <=32'hFF22001E;14'd16082:data <=32'hFF370044;
14'd16083:data <=32'hFF580062;14'd16084:data <=32'hFF7C0075;14'd16085:data <=32'hFFA0007D;
14'd16086:data <=32'hFFC2007A;14'd16087:data <=32'hFFDD006D;14'd16088:data <=32'hFFEF005D;
14'd16089:data <=32'hFFFB004E;14'd16090:data <=32'h00010040;14'd16091:data <=32'h00030035;
14'd16092:data <=32'h0007002C;14'd16093:data <=32'h00080022;14'd16094:data <=32'h000A0018;
14'd16095:data <=32'h0009000B;14'd16096:data <=32'h0003FFFF;14'd16097:data <=32'hFFF8FFF3;
14'd16098:data <=32'hFFE9FFEB;14'd16099:data <=32'hFFD6FFEA;14'd16100:data <=32'hFFC3FFEF;
14'd16101:data <=32'hFFB2FFFB;14'd16102:data <=32'hFFA4000B;14'd16103:data <=32'hFF9A0021;
14'd16104:data <=32'hFF960038;14'd16105:data <=32'hFF97004F;14'd16106:data <=32'hFF9E0069;
14'd16107:data <=32'hFFAA0081;14'd16108:data <=32'hFFBD0099;14'd16109:data <=32'hFFD600AF;
14'd16110:data <=32'hFFF600BE;14'd16111:data <=32'h001D00C4;14'd16112:data <=32'h004600C0;
14'd16113:data <=32'h006E00AF;14'd16114:data <=32'h008C0093;14'd16115:data <=32'h00A10070;
14'd16116:data <=32'h00AA004A;14'd16117:data <=32'h00A70026;14'd16118:data <=32'h009B0009;
14'd16119:data <=32'h0089FFF5;14'd16120:data <=32'h0076FFEB;14'd16121:data <=32'h0065FFE7;
14'd16122:data <=32'h0058FFE9;14'd16123:data <=32'h0050FFED;14'd16124:data <=32'h004CFFF3;
14'd16125:data <=32'h004DFFF9;14'd16126:data <=32'h0052FFFF;14'd16127:data <=32'h005C0004;
14'd16128:data <=32'h007CFFFA;14'd16129:data <=32'h0091FFEE;14'd16130:data <=32'h0090FFDC;
14'd16131:data <=32'h005FFFD8;14'd16132:data <=32'h00A2FFC3;14'd16133:data <=32'h00A0FFA4;
14'd16134:data <=32'h0094FF83;14'd16135:data <=32'h007FFF67;14'd16136:data <=32'h0061FF51;
14'd16137:data <=32'h0040FF46;14'd16138:data <=32'h001FFF44;14'd16139:data <=32'h0002FF49;
14'd16140:data <=32'hFFEAFF53;14'd16141:data <=32'hFFD6FF5E;14'd16142:data <=32'hFFC6FF6A;
14'd16143:data <=32'hFFB7FF76;14'd16144:data <=32'hFFA9FF83;14'd16145:data <=32'hFF9DFF92;
14'd16146:data <=32'hFF95FFA4;14'd16147:data <=32'hFF90FFB6;14'd16148:data <=32'hFF8EFFC6;
14'd16149:data <=32'hFF90FFD5;14'd16150:data <=32'hFF92FFE0;14'd16151:data <=32'hFF93FFE9;
14'd16152:data <=32'hFF93FFF3;14'd16153:data <=32'hFF92FFFF;14'd16154:data <=32'hFF93000D;
14'd16155:data <=32'hFF97001F;14'd16156:data <=32'hFFA20030;14'd16157:data <=32'hFFB3003F;
14'd16158:data <=32'hFFCB0046;14'd16159:data <=32'hFFE30045;14'd16160:data <=32'hFFF9003A;
14'd16161:data <=32'h000A0029;14'd16162:data <=32'h00120013;14'd16163:data <=32'h0012FFFB;
14'd16164:data <=32'h0007FFE6;14'd16165:data <=32'hFFF7FFD5;14'd16166:data <=32'hFFE2FFCB;
14'd16167:data <=32'hFFCBFFC7;14'd16168:data <=32'hFFB1FFCB;14'd16169:data <=32'hFF98FFD5;
14'd16170:data <=32'hFF82FFE7;14'd16171:data <=32'hFF700000;14'd16172:data <=32'hFF63001F;
14'd16173:data <=32'hFF5E0043;14'd16174:data <=32'hFF65006A;14'd16175:data <=32'hFF78008E;
14'd16176:data <=32'hFF9300AC;14'd16177:data <=32'hFFB700C0;14'd16178:data <=32'hFFDE00CA;
14'd16179:data <=32'h000300C8;14'd16180:data <=32'h002300BE;14'd16181:data <=32'h003B00AD;
14'd16182:data <=32'h004D009C;14'd16183:data <=32'h0059008D;14'd16184:data <=32'h00630080;
14'd16185:data <=32'h006B0075;14'd16186:data <=32'h0075006B;14'd16187:data <=32'h007F0060;
14'd16188:data <=32'h00890053;14'd16189:data <=32'h00920044;14'd16190:data <=32'h00990035;
14'd16191:data <=32'h009D0027;14'd16192:data <=32'h00140021;14'd16193:data <=32'h0027003E;
14'd16194:data <=32'h004A0045;14'd16195:data <=32'h00AAFFF2;14'd16196:data <=32'h00E1FFD3;
14'd16197:data <=32'h00D4FFAC;14'd16198:data <=32'h00BCFF89;14'd16199:data <=32'h009DFF6C;
14'd16200:data <=32'h0075FF5B;14'd16201:data <=32'h004DFF56;14'd16202:data <=32'h0028FF5F;
14'd16203:data <=32'h000AFF70;14'd16204:data <=32'hFFF9FF87;14'd16205:data <=32'hFFF1FF9C;
14'd16206:data <=32'hFFF1FFAE;14'd16207:data <=32'hFFF7FFBB;14'd16208:data <=32'hFFFEFFC2;
14'd16209:data <=32'h0003FFC5;14'd16210:data <=32'h0009FFC3;14'd16211:data <=32'h000DFFBE;
14'd16212:data <=32'h000FFFB7;14'd16213:data <=32'h000EFFAE;14'd16214:data <=32'h0009FFA2;
14'd16215:data <=32'hFFFEFF97;14'd16216:data <=32'hFFECFF8D;14'd16217:data <=32'hFFD6FF8B;
14'd16218:data <=32'hFFBDFF90;14'd16219:data <=32'hFFA6FF9E;14'd16220:data <=32'hFF95FFB5;
14'd16221:data <=32'hFF8DFFD0;14'd16222:data <=32'hFF8FFFEC;14'd16223:data <=32'hFF9A0004;
14'd16224:data <=32'hFFAC0013;14'd16225:data <=32'hFFBF001C;14'd16226:data <=32'hFFD3001B;
14'd16227:data <=32'hFFE20016;14'd16228:data <=32'hFFEC000C;14'd16229:data <=32'hFFF20000;
14'd16230:data <=32'hFFF4FFF5;14'd16231:data <=32'hFFF1FFE9;14'd16232:data <=32'hFFEDFFDE;
14'd16233:data <=32'hFFE3FFD4;14'd16234:data <=32'hFFD6FFCB;14'd16235:data <=32'hFFC6FFC8;
14'd16236:data <=32'hFFB2FFC8;14'd16237:data <=32'hFF9FFFCF;14'd16238:data <=32'hFF8DFFDC;
14'd16239:data <=32'hFF7FFFEF;14'd16240:data <=32'hFF770004;14'd16241:data <=32'hFF740019;
14'd16242:data <=32'hFF75002D;14'd16243:data <=32'hFF78003E;14'd16244:data <=32'hFF7B004E;
14'd16245:data <=32'hFF7C005E;14'd16246:data <=32'hFF7F0072;14'd16247:data <=32'hFF840088;
14'd16248:data <=32'hFF8D00A4;14'd16249:data <=32'hFF9F00C2;14'd16250:data <=32'hFFBB00DE;
14'd16251:data <=32'hFFE000F4;14'd16252:data <=32'h000C0100;14'd16253:data <=32'h003B0102;
14'd16254:data <=32'h006A00F9;14'd16255:data <=32'h009600E6;14'd16256:data <=32'h00220026;
14'd16257:data <=32'h001E003F;14'd16258:data <=32'h002F006A;14'd16259:data <=32'h00BC00B6;
14'd16260:data <=32'h01150089;14'd16261:data <=32'h0124004C;14'd16262:data <=32'h0124000E;
14'd16263:data <=32'h0113FFD4;14'd16264:data <=32'h00F3FFA1;14'd16265:data <=32'h00C6FF7D;
14'd16266:data <=32'h0096FF69;14'd16267:data <=32'h0069FF66;14'd16268:data <=32'h0041FF6F;
14'd16269:data <=32'h0024FF80;14'd16270:data <=32'h0011FF94;14'd16271:data <=32'h0007FFA7;
14'd16272:data <=32'h0004FFB9;14'd16273:data <=32'h0004FFC7;14'd16274:data <=32'h0007FFD1;
14'd16275:data <=32'h000DFFDA;14'd16276:data <=32'h0016FFDF;14'd16277:data <=32'h0020FFDF;
14'd16278:data <=32'h002AFFD9;14'd16279:data <=32'h002FFFCE;14'd16280:data <=32'h0030FFC0;
14'd16281:data <=32'h002AFFB1;14'd16282:data <=32'h001EFFA6;14'd16283:data <=32'h000EFF9F;
14'd16284:data <=32'hFFFDFFA0;14'd16285:data <=32'hFFEFFFA6;14'd16286:data <=32'hFFE5FFAE;
14'd16287:data <=32'hFFE0FFB8;14'd16288:data <=32'hFFDFFFC0;14'd16289:data <=32'hFFE0FFC5;
14'd16290:data <=32'hFFE1FFC6;14'd16291:data <=32'hFFDFFFC5;14'd16292:data <=32'hFFDAFFC6;
14'd16293:data <=32'hFFD4FFC7;14'd16294:data <=32'hFFCDFFCB;14'd16295:data <=32'hFFC9FFD2;
14'd16296:data <=32'hFFC7FFDA;14'd16297:data <=32'hFFC9FFE1;14'd16298:data <=32'hFFCCFFE6;
14'd16299:data <=32'hFFD0FFE7;14'd16300:data <=32'hFFD3FFE8;14'd16301:data <=32'hFFD6FFE5;
14'd16302:data <=32'hFFD6FFE2;14'd16303:data <=32'hFFD4FFDE;14'd16304:data <=32'hFFD3FFDA;
14'd16305:data <=32'hFFCFFFD3;14'd16306:data <=32'hFFC9FFCB;14'd16307:data <=32'hFFBDFFC2;
14'd16308:data <=32'hFFABFFB9;14'd16309:data <=32'hFF91FFB6;14'd16310:data <=32'hFF71FFBB;
14'd16311:data <=32'hFF4EFFCC;14'd16312:data <=32'hFF2EFFEB;14'd16313:data <=32'hFF170016;
14'd16314:data <=32'hFF0C004B;14'd16315:data <=32'hFF100083;14'd16316:data <=32'hFF2500BA;
14'd16317:data <=32'hFF4800EA;14'd16318:data <=32'hFF760111;14'd16319:data <=32'hFFAC012C;
14'd16320:data <=32'hFFDB0090;14'd16321:data <=32'hFFE200AD;14'd16322:data <=32'hFFE000CC;
14'd16323:data <=32'hFFDA011A;14'd16324:data <=32'h004C0119;14'd16325:data <=32'h007E00FF;
14'd16326:data <=32'h00A500DB;14'd16327:data <=32'h00C300B0;14'd16328:data <=32'h00D20081;
14'd16329:data <=32'h00D20054;14'd16330:data <=32'h00CA002E;14'd16331:data <=32'h00BB0012;
14'd16332:data <=32'h00ABFFFD;14'd16333:data <=32'h009EFFEE;14'd16334:data <=32'h0092FFE2;
14'd16335:data <=32'h0088FFD6;14'd16336:data <=32'h007DFFCB;14'd16337:data <=32'h0071FFBF;
14'd16338:data <=32'h0062FFB6;14'd16339:data <=32'h0052FFAF;14'd16340:data <=32'h0042FFAE;
14'd16341:data <=32'h0033FFB0;14'd16342:data <=32'h0028FFB4;14'd16343:data <=32'h001FFFB9;
14'd16344:data <=32'h0018FFBD;14'd16345:data <=32'h0010FFC1;14'd16346:data <=32'h000AFFC6;
14'd16347:data <=32'h0004FFCE;14'd16348:data <=32'h0001FFD8;14'd16349:data <=32'h0002FFE3;
14'd16350:data <=32'h0007FFEE;14'd16351:data <=32'h0014FFF5;14'd16352:data <=32'h0023FFF6;
14'd16353:data <=32'h0032FFEE;14'd16354:data <=32'h003DFFDF;14'd16355:data <=32'h0042FFCB;
14'd16356:data <=32'h003FFFB7;14'd16357:data <=32'h0033FFA4;14'd16358:data <=32'h0022FF97;
14'd16359:data <=32'h000EFF90;14'd16360:data <=32'hFFF9FF90;14'd16361:data <=32'hFFE7FF95;
14'd16362:data <=32'hFFD9FF9F;14'd16363:data <=32'hFFD0FFA9;14'd16364:data <=32'hFFCAFFB5;
14'd16365:data <=32'hFFC7FFC0;14'd16366:data <=32'hFFC7FFCA;14'd16367:data <=32'hFFCBFFD2;
14'd16368:data <=32'hFFD0FFD8;14'd16369:data <=32'hFFD9FFD9;14'd16370:data <=32'hFFE1FFD5;
14'd16371:data <=32'hFFE6FFCA;14'd16372:data <=32'hFFE5FFBA;14'd16373:data <=32'hFFDBFFA7;
14'd16374:data <=32'hFFC7FF97;14'd16375:data <=32'hFFAAFF8C;14'd16376:data <=32'hFF87FF8E;
14'd16377:data <=32'hFF62FF9C;14'd16378:data <=32'hFF41FFB6;14'd16379:data <=32'hFF28FFDB;
14'd16380:data <=32'hFF1B0005;14'd16381:data <=32'hFF190030;14'd16382:data <=32'hFF21005B;
14'd16383:data <=32'hFF320081;
        
        endcase
        
end    
    
    assign dout = data;
    
endmodule
