`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 05/23/2023 02:45:31 PM
// Design Name: 
// Module Name: rom
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module sp_rom #(
    parameter integer ADDRW = 14,
    parameter integer DATA_WIDTH = 32,
    parameter RAM_TYPE = "block"
)
(
input [ADDRW-1:0] addr,
input clk,
input en,
output wire [DATA_WIDTH-1:0] dout
    );
    
//DD clock
//(*ram_style = "registers"*)reg r_clk50=0;

//wire w_xor_clk50=(r_clk50 ^ clk);

//always@(posedge w_xor_clk50) begin

//    r_clk50=~r_clk50;

//    // your code on both neg/pos
//end
 
    
 (*rom_style = RAM_TYPE*) reg [DATA_WIDTH-1:0] data;   
    
always@(negedge clk)
begin
    if(en)
    case (addr)
    14'd0:data <=32'h00000000;14'd1:data <=32'hFFF1FFD0;14'd2:data <=32'hFFE1FFAE;
14'd3:data <=32'hFFDFFFA6;14'd4:data <=32'hFFC4FFB3;14'd5:data <=32'hFFBBFFBF;
14'd6:data <=32'hFFB5FFCB;14'd7:data <=32'hFFAFFFD8;14'd8:data <=32'hFFAFFFE5;
14'd9:data <=32'hFFB0FFEF;14'd10:data <=32'hFFB3FFF7;14'd11:data <=32'hFFB4FFFD;
14'd12:data <=32'hFFB40004;14'd13:data <=32'hFFB3000C;14'd14:data <=32'hFFB40015;
14'd15:data <=32'hFFB60021;14'd16:data <=32'hFFBB002D;14'd17:data <=32'hFFC40037;
14'd18:data <=32'hFFCF003F;14'd19:data <=32'hFFDC0044;14'd20:data <=32'hFFE90046;
14'd21:data <=32'hFFF60045;14'd22:data <=32'h00010041;14'd23:data <=32'h000B003B;
14'd24:data <=32'h00140035;14'd25:data <=32'h001B002B;14'd26:data <=32'h00200020;
14'd27:data <=32'h00210015;14'd28:data <=32'h001F0009;14'd29:data <=32'h0018FFFE;
14'd30:data <=32'h000EFFF7;14'd31:data <=32'h0002FFF5;14'd32:data <=32'hFFF6FFF8;
14'd33:data <=32'hFFECFFFF;14'd34:data <=32'hFFE70009;14'd35:data <=32'hFFE50015;
14'd36:data <=32'hFFE80020;14'd37:data <=32'hFFEF0029;14'd38:data <=32'hFFF7002F;
14'd39:data <=32'h00000032;14'd40:data <=32'h00090033;14'd41:data <=32'h00120032;
14'd42:data <=32'h0019002F;14'd43:data <=32'h0020002B;14'd44:data <=32'h00260026;
14'd45:data <=32'h002A0021;14'd46:data <=32'h002D001B;14'd47:data <=32'h002F0014;
14'd48:data <=32'h002F000F;14'd49:data <=32'h002E000B;14'd50:data <=32'h002C0009;
14'd51:data <=32'h002D0008;14'd52:data <=32'h002F0008;14'd53:data <=32'h00330007;
14'd54:data <=32'h00390004;14'd55:data <=32'h003FFFFE;14'd56:data <=32'h0044FFF4;
14'd57:data <=32'h0047FFE8;14'd58:data <=32'h0045FFDB;14'd59:data <=32'h003FFFCE;
14'd60:data <=32'h0037FFC4;14'd61:data <=32'h002DFFBD;14'd62:data <=32'h0022FFB8;
14'd63:data <=32'h0018FFB6;14'd64:data <=32'h005DFFC2;14'd65:data <=32'h0056FFA4;
14'd66:data <=32'h0044FF91;14'd67:data <=32'h0014FFBB;14'd68:data <=32'hFFFAFFCE;
14'd69:data <=32'hFFF8FFD1;14'd70:data <=32'hFFF8FFD4;14'd71:data <=32'hFFF9FFD5;
14'd72:data <=32'hFFFAFFD3;14'd73:data <=32'hFFFAFFCF;14'd74:data <=32'hFFF8FFC9;
14'd75:data <=32'hFFF2FFC2;14'd76:data <=32'hFFE7FFBC;14'd77:data <=32'hFFD9FFBA;
14'd78:data <=32'hFFC8FFBD;14'd79:data <=32'hFFB8FFC6;14'd80:data <=32'hFFABFFD4;
14'd81:data <=32'hFFA2FFE5;14'd82:data <=32'hFF9FFFF8;14'd83:data <=32'hFFA2000B;
14'd84:data <=32'hFFA8001C;14'd85:data <=32'hFFB1002B;14'd86:data <=32'hFFBD0037;
14'd87:data <=32'hFFCC003F;14'd88:data <=32'hFFDB0045;14'd89:data <=32'hFFEC0046;
14'd90:data <=32'hFFFC0042;14'd91:data <=32'h000A003B;14'd92:data <=32'h0016002E;
14'd93:data <=32'h001C0020;14'd94:data <=32'h001C0012;14'd95:data <=32'h00180005;
14'd96:data <=32'h0010FFFB;14'd97:data <=32'h0006FFF6;14'd98:data <=32'hFFFCFFF5;
14'd99:data <=32'hFFF3FFF7;14'd100:data <=32'hFFECFFFB;14'd101:data <=32'hFFE70000;
14'd102:data <=32'hFFE40006;14'd103:data <=32'hFFE1000B;14'd104:data <=32'hFFDF0012;
14'd105:data <=32'hFFDE0018;14'd106:data <=32'hFFDE0020;14'd107:data <=32'hFFDF0029;
14'd108:data <=32'hFFE30033;14'd109:data <=32'hFFE9003B;14'd110:data <=32'hFFF20042;
14'd111:data <=32'hFFFD0048;14'd112:data <=32'h0008004B;14'd113:data <=32'h0014004D;
14'd114:data <=32'h0020004C;14'd115:data <=32'h002D004A;14'd116:data <=32'h003A0046;
14'd117:data <=32'h0048003F;14'd118:data <=32'h00550035;14'd119:data <=32'h00600026;
14'd120:data <=32'h00690014;14'd121:data <=32'h006CFFFF;14'd122:data <=32'h0069FFEA;
14'd123:data <=32'h0060FFD6;14'd124:data <=32'h0053FFC6;14'd125:data <=32'h0043FFBC;
14'd126:data <=32'h0031FFB7;14'd127:data <=32'h0022FFB8;14'd128:data <=32'h00550009;
14'd129:data <=32'h0063FFF4;14'd130:data <=32'h0062FFD7;14'd131:data <=32'h0021FFBA;
14'd132:data <=32'h0003FFD0;14'd133:data <=32'h0000FFD8;14'd134:data <=32'h0001FFDF;
14'd135:data <=32'h0004FFE4;14'd136:data <=32'h000AFFE7;14'd137:data <=32'h0010FFE6;
14'd138:data <=32'h0016FFE0;14'd139:data <=32'h0019FFD7;14'd140:data <=32'h0017FFCC;
14'd141:data <=32'h0010FFC1;14'd142:data <=32'h0004FFB8;14'd143:data <=32'hFFF6FFB4;
14'd144:data <=32'hFFE6FFB5;14'd145:data <=32'hFFD8FFBB;14'd146:data <=32'hFFCCFFC4;
14'd147:data <=32'hFFC4FFCF;14'd148:data <=32'hFFBEFFDA;14'd149:data <=32'hFFBBFFE6;
14'd150:data <=32'hFFBAFFF2;14'd151:data <=32'hFFBBFFFD;14'd152:data <=32'hFFBE0009;
14'd153:data <=32'hFFC40013;14'd154:data <=32'hFFCD001B;14'd155:data <=32'hFFD60021;
14'd156:data <=32'hFFE10023;14'd157:data <=32'hFFEB0022;14'd158:data <=32'hFFF2001F;
14'd159:data <=32'hFFF8001A;14'd160:data <=32'hFFFB0015;14'd161:data <=32'hFFFC0011;
14'd162:data <=32'hFFFD000E;14'd163:data <=32'hFFFE000B;14'd164:data <=32'hFFFF0008;
14'd165:data <=32'hFFFF0003;14'd166:data <=32'hFFFFFFFE;14'd167:data <=32'hFFFCFFF9;
14'd168:data <=32'hFFF7FFF3;14'd169:data <=32'hFFEEFFEF;14'd170:data <=32'hFFE4FFED;
14'd171:data <=32'hFFD7FFF0;14'd172:data <=32'hFFCCFFF8;14'd173:data <=32'hFFC30002;
14'd174:data <=32'hFFBC0011;14'd175:data <=32'hFFBA0021;14'd176:data <=32'hFFBB0032;
14'd177:data <=32'hFFC10043;14'd178:data <=32'hFFCB0054;14'd179:data <=32'hFFD90062;
14'd180:data <=32'hFFEB006E;14'd181:data <=32'h00000076;14'd182:data <=32'h00190079;
14'd183:data <=32'h00330075;14'd184:data <=32'h004B006A;14'd185:data <=32'h00610059;
14'd186:data <=32'h00700042;14'd187:data <=32'h00770028;14'd188:data <=32'h0078000F;
14'd189:data <=32'h0072FFF8;14'd190:data <=32'h0067FFE6;14'd191:data <=32'h005AFFD8;
14'd192:data <=32'h0040000D;14'd193:data <=32'h004A0005;14'd194:data <=32'h0056FFF7;
14'd195:data <=32'h0060FFD6;14'd196:data <=32'h0041FFDE;14'd197:data <=32'h003AFFD9;
14'd198:data <=32'h0033FFD6;14'd199:data <=32'h002DFFD5;14'd200:data <=32'h0029FFD3;
14'd201:data <=32'h0026FFD2;14'd202:data <=32'h0023FFD0;14'd203:data <=32'h0020FFCC;
14'd204:data <=32'h001CFFC6;14'd205:data <=32'h0014FFC1;14'd206:data <=32'h000BFFBE;
14'd207:data <=32'hFFFFFFBE;14'd208:data <=32'hFFF4FFC1;14'd209:data <=32'hFFEBFFC8;
14'd210:data <=32'hFFE5FFD0;14'd211:data <=32'hFFE3FFD8;14'd212:data <=32'hFFE3FFE0;
14'd213:data <=32'hFFE4FFE5;14'd214:data <=32'hFFE6FFE9;14'd215:data <=32'hFFE8FFEA;
14'd216:data <=32'hFFE8FFEC;14'd217:data <=32'hFFE8FFED;14'd218:data <=32'hFFE8FFEE;
14'd219:data <=32'hFFE8FFF0;14'd220:data <=32'hFFE8FFF0;14'd221:data <=32'hFFE8FFF1;
14'd222:data <=32'hFFE6FFF1;14'd223:data <=32'hFFE4FFF2;14'd224:data <=32'hFFE1FFF4;
14'd225:data <=32'hFFDEFFF8;14'd226:data <=32'hFFDDFFFE;14'd227:data <=32'hFFDF0004;
14'd228:data <=32'hFFE3000A;14'd229:data <=32'hFFE9000D;14'd230:data <=32'hFFF1000E;
14'd231:data <=32'hFFF8000B;14'd232:data <=32'hFFFD0004;14'd233:data <=32'hFFFFFFFB;
14'd234:data <=32'hFFFCFFF2;14'd235:data <=32'hFFF5FFEA;14'd236:data <=32'hFFEBFFE5;
14'd237:data <=32'hFFE0FFE4;14'd238:data <=32'hFFD4FFE7;14'd239:data <=32'hFFC9FFED;
14'd240:data <=32'hFFBFFFF6;14'd241:data <=32'hFFB70002;14'd242:data <=32'hFFB10010;
14'd243:data <=32'hFFB00020;14'd244:data <=32'hFFB10032;14'd245:data <=32'hFFB70044;
14'd246:data <=32'hFFC30054;14'd247:data <=32'hFFD30062;14'd248:data <=32'hFFE6006B;
14'd249:data <=32'hFFFB006E;14'd250:data <=32'h000F006C;14'd251:data <=32'h00210065;
14'd252:data <=32'h002F005B;14'd253:data <=32'h003A0050;14'd254:data <=32'h00400045;
14'd255:data <=32'h0045003B;14'd256:data <=32'h0051002D;14'd257:data <=32'h00590023;
14'd258:data <=32'h005E001E;14'd259:data <=32'h00590040;14'd260:data <=32'h004F0043;
14'd261:data <=32'h005A0037;14'd262:data <=32'h00630029;14'd263:data <=32'h006A0018;
14'd264:data <=32'h006D0007;14'd265:data <=32'h006DFFF5;14'd266:data <=32'h006AFFE3;
14'd267:data <=32'h0064FFD1;14'd268:data <=32'h0059FFC0;14'd269:data <=32'h004AFFB1;
14'd270:data <=32'h0036FFA6;14'd271:data <=32'h0020FFA1;14'd272:data <=32'h000AFFA3;
14'd273:data <=32'hFFF7FFAB;14'd274:data <=32'hFFE7FFB8;14'd275:data <=32'hFFDFFFC8;
14'd276:data <=32'hFFDBFFD8;14'd277:data <=32'hFFDDFFE6;14'd278:data <=32'hFFE2FFF1;
14'd279:data <=32'hFFE9FFF8;14'd280:data <=32'hFFF0FFFD;14'd281:data <=32'hFFF8FFFF;
14'd282:data <=32'hFFFEFFFF;14'd283:data <=32'h0005FFFC;14'd284:data <=32'h000AFFF7;
14'd285:data <=32'h000CFFF1;14'd286:data <=32'h000DFFEA;14'd287:data <=32'h000BFFE3;
14'd288:data <=32'h0005FFDD;14'd289:data <=32'hFFFEFFD9;14'd290:data <=32'hFFF6FFD9;
14'd291:data <=32'hFFEFFFDB;14'd292:data <=32'hFFE9FFE0;14'd293:data <=32'hFFE7FFE6;
14'd294:data <=32'hFFE7FFEA;14'd295:data <=32'hFFE8FFEE;14'd296:data <=32'hFFEAFFEF;
14'd297:data <=32'hFFECFFED;14'd298:data <=32'hFFEBFFEB;14'd299:data <=32'hFFE9FFE9;
14'd300:data <=32'hFFE4FFE8;14'd301:data <=32'hFFDFFFE9;14'd302:data <=32'hFFDAFFEA;
14'd303:data <=32'hFFD5FFEE;14'd304:data <=32'hFFD2FFF3;14'd305:data <=32'hFFCFFFF7;
14'd306:data <=32'hFFCCFFFC;14'd307:data <=32'hFFCA0002;14'd308:data <=32'hFFC80007;
14'd309:data <=32'hFFC7000F;14'd310:data <=32'hFFC70016;14'd311:data <=32'hFFC9001E;
14'd312:data <=32'hFFCD0024;14'd313:data <=32'hFFD2002A;14'd314:data <=32'hFFD7002D;
14'd315:data <=32'hFFDA0030;14'd316:data <=32'hFFDC0032;14'd317:data <=32'hFFDD0036;
14'd318:data <=32'hFFDD003D;14'd319:data <=32'hFFDF0046;14'd320:data <=32'h00140063;
14'd321:data <=32'h00240063;14'd322:data <=32'h002A005D;14'd323:data <=32'hFFF5005B;
14'd324:data <=32'hFFEF0071;14'd325:data <=32'h00050078;14'd326:data <=32'h001C0079;
14'd327:data <=32'h00340073;14'd328:data <=32'h0049006A;14'd329:data <=32'h005D005B;
14'd330:data <=32'h006E0048;14'd331:data <=32'h007A0032;14'd332:data <=32'h00810017;
14'd333:data <=32'h0080FFFC;14'd334:data <=32'h0079FFE2;14'd335:data <=32'h006AFFCB;
14'd336:data <=32'h0056FFBB;14'd337:data <=32'h003FFFB1;14'd338:data <=32'h0029FFAF;
14'd339:data <=32'h0015FFB3;14'd340:data <=32'h0006FFBB;14'd341:data <=32'hFFFBFFC5;
14'd342:data <=32'hFFF3FFCF;14'd343:data <=32'hFFEFFFDA;14'd344:data <=32'hFFEEFFE3;
14'd345:data <=32'hFFEEFFEC;14'd346:data <=32'hFFF0FFF4;14'd347:data <=32'hFFF4FFFB;
14'd348:data <=32'hFFF90000;14'd349:data <=32'h00000003;14'd350:data <=32'h00080003;
14'd351:data <=32'h000E0001;14'd352:data <=32'h0013FFFD;14'd353:data <=32'h0016FFF7;
14'd354:data <=32'h0018FFF2;14'd355:data <=32'h0018FFED;14'd356:data <=32'h0017FFE9;
14'd357:data <=32'h0016FFE4;14'd358:data <=32'h0016FFDF;14'd359:data <=32'h0015FFDA;
14'd360:data <=32'h0012FFD3;14'd361:data <=32'h000DFFCB;14'd362:data <=32'h0006FFC5;
14'd363:data <=32'hFFFBFFBF;14'd364:data <=32'hFFEEFFBD;14'd365:data <=32'hFFE1FFBF;
14'd366:data <=32'hFFD3FFC5;14'd367:data <=32'hFFCAFFCE;14'd368:data <=32'hFFC2FFD9;
14'd369:data <=32'hFFBFFFE5;14'd370:data <=32'hFFBEFFF1;14'd371:data <=32'hFFC1FFFB;
14'd372:data <=32'hFFC40004;14'd373:data <=32'hFFCA000A;14'd374:data <=32'hFFCF000F;
14'd375:data <=32'hFFD60013;14'd376:data <=32'hFFDC0013;14'd377:data <=32'hFFE20011;
14'd378:data <=32'hFFE5000D;14'd379:data <=32'hFFE50007;14'd380:data <=32'hFFE20002;
14'd381:data <=32'hFFD9FFFF;14'd382:data <=32'hFFCEFFFF;14'd383:data <=32'hFFC30006;
14'd384:data <=32'hFFC4002F;14'd385:data <=32'hFFC4003D;14'd386:data <=32'hFFCC0042;
14'd387:data <=32'hFFCD0025;14'd388:data <=32'hFFBA003F;14'd389:data <=32'hFFC4004E;
14'd390:data <=32'hFFD1005A;14'd391:data <=32'hFFE10062;14'd392:data <=32'hFFF30068;
14'd393:data <=32'h0004006A;14'd394:data <=32'h00170068;14'd395:data <=32'h00290062;
14'd396:data <=32'h003A0058;14'd397:data <=32'h0048004A;14'd398:data <=32'h00510038;
14'd399:data <=32'h00550027;14'd400:data <=32'h00540015;14'd401:data <=32'h00500007;
14'd402:data <=32'h0049FFFC;14'd403:data <=32'h0041FFF4;14'd404:data <=32'h003BFFF0;
14'd405:data <=32'h0035FFEB;14'd406:data <=32'h0030FFE7;14'd407:data <=32'h002BFFE3;
14'd408:data <=32'h0025FFDF;14'd409:data <=32'h001DFFDC;14'd410:data <=32'h0015FFDB;
14'd411:data <=32'h000CFFDC;14'd412:data <=32'h0004FFE0;14'd413:data <=32'hFFFFFFE5;
14'd414:data <=32'hFFFBFFED;14'd415:data <=32'hFFFAFFF4;14'd416:data <=32'hFFFAFFFA;
14'd417:data <=32'hFFFD0000;14'd418:data <=32'h00010006;14'd419:data <=32'h0006000A;
14'd420:data <=32'h000D000E;14'd421:data <=32'h0016000F;14'd422:data <=32'h0021000E;
14'd423:data <=32'h002C0008;14'd424:data <=32'h0035FFFE;14'd425:data <=32'h003CFFF0;
14'd426:data <=32'h003EFFE0;14'd427:data <=32'h003BFFCF;14'd428:data <=32'h0031FFBF;
14'd429:data <=32'h0024FFB2;14'd430:data <=32'h0013FFAB;14'd431:data <=32'h0002FFA8;
14'd432:data <=32'hFFF1FFAA;14'd433:data <=32'hFFE2FFB0;14'd434:data <=32'hFFD6FFB8;
14'd435:data <=32'hFFCDFFC2;14'd436:data <=32'hFFC7FFCD;14'd437:data <=32'hFFC3FFD7;
14'd438:data <=32'hFFC2FFE2;14'd439:data <=32'hFFC2FFEC;14'd440:data <=32'hFFC5FFF4;
14'd441:data <=32'hFFCAFFFA;14'd442:data <=32'hFFCFFFFE;14'd443:data <=32'hFFD4FFFE;
14'd444:data <=32'hFFD6FFFC;14'd445:data <=32'hFFD4FFF9;14'd446:data <=32'hFFCFFFF8;
14'd447:data <=32'hFFC8FFF9;14'd448:data <=32'hFFDDFFE5;14'd449:data <=32'hFFCBFFE6;
14'd450:data <=32'hFFC0FFF2;14'd451:data <=32'hFFCA001A;14'd452:data <=32'hFFB8002F;
14'd453:data <=32'hFFC20039;14'd454:data <=32'hFFCE0040;14'd455:data <=32'hFFDA0043;
14'd456:data <=32'hFFE50044;14'd457:data <=32'hFFEE0043;14'd458:data <=32'hFFF60041;
14'd459:data <=32'hFFFE003F;14'd460:data <=32'h0005003B;14'd461:data <=32'h000A0036;
14'd462:data <=32'h000F0031;14'd463:data <=32'h0011002C;14'd464:data <=32'h00110028;
14'd465:data <=32'h000F0026;14'd466:data <=32'h000E0026;14'd467:data <=32'h000F0029;
14'd468:data <=32'h0013002C;14'd469:data <=32'h001A002E;14'd470:data <=32'h0023002D;
14'd471:data <=32'h002D0028;14'd472:data <=32'h00350020;14'd473:data <=32'h003A0015;
14'd474:data <=32'h003B0009;14'd475:data <=32'h0039FFFD;14'd476:data <=32'h0033FFF3;
14'd477:data <=32'h002CFFEC;14'd478:data <=32'h0023FFE7;14'd479:data <=32'h001AFFE5;
14'd480:data <=32'h0011FFE6;14'd481:data <=32'h0009FFE8;14'd482:data <=32'h0001FFEE;
14'd483:data <=32'hFFFCFFF5;14'd484:data <=32'hFFF9FFFE;14'd485:data <=32'hFFFB0008;
14'd486:data <=32'h00000012;14'd487:data <=32'h00090019;14'd488:data <=32'h0015001D;
14'd489:data <=32'h0022001C;14'd490:data <=32'h002E0016;14'd491:data <=32'h0038000C;
14'd492:data <=32'h003F0000;14'd493:data <=32'h0041FFF3;14'd494:data <=32'h0040FFE6;
14'd495:data <=32'h003CFFDB;14'd496:data <=32'h0036FFD2;14'd497:data <=32'h0030FFCB;
14'd498:data <=32'h002AFFC4;14'd499:data <=32'h0022FFBE;14'd500:data <=32'h001BFFB8;
14'd501:data <=32'h0012FFB3;14'd502:data <=32'h0007FFAF;14'd503:data <=32'hFFFCFFAD;
14'd504:data <=32'hFFF1FFAC;14'd505:data <=32'hFFE5FFAE;14'd506:data <=32'hFFDBFFB1;
14'd507:data <=32'hFFD1FFB5;14'd508:data <=32'hFFC6FFB9;14'd509:data <=32'hFFBCFFBF;
14'd510:data <=32'hFFB1FFC7;14'd511:data <=32'hFFA6FFD2;14'd512:data <=32'hFFFEFFE8;
14'd513:data <=32'hFFF3FFDA;14'd514:data <=32'hFFDEFFD4;14'd515:data <=32'hFF9CFFF5;
14'd516:data <=32'hFF880015;14'd517:data <=32'hFF95002B;14'd518:data <=32'hFFA5003B;
14'd519:data <=32'hFFB90045;14'd520:data <=32'hFFCC0049;14'd521:data <=32'hFFDD0049;
14'd522:data <=32'hFFEC0044;14'd523:data <=32'hFFF7003E;14'd524:data <=32'h00010036;
14'd525:data <=32'h0007002C;14'd526:data <=32'h00090022;14'd527:data <=32'h00080018;
14'd528:data <=32'h00030011;14'd529:data <=32'hFFFC000D;14'd530:data <=32'hFFF4000D;
14'd531:data <=32'hFFED0012;14'd532:data <=32'hFFE9001A;14'd533:data <=32'hFFE90024;
14'd534:data <=32'hFFEE002D;14'd535:data <=32'hFFF70034;14'd536:data <=32'h00020037;
14'd537:data <=32'h000C0036;14'd538:data <=32'h00160032;14'd539:data <=32'h001D002C;
14'd540:data <=32'h00220025;14'd541:data <=32'h0024001E;14'd542:data <=32'h00260017;
14'd543:data <=32'h00260011;14'd544:data <=32'h0025000B;14'd545:data <=32'h00220005;
14'd546:data <=32'h001F0000;14'd547:data <=32'h0019FFFD;14'd548:data <=32'h0014FFFC;
14'd549:data <=32'h000FFFFE;14'd550:data <=32'h000B0001;14'd551:data <=32'h000A0005;
14'd552:data <=32'h000A000A;14'd553:data <=32'h000D000E;14'd554:data <=32'h00110010;
14'd555:data <=32'h00140010;14'd556:data <=32'h0018000F;14'd557:data <=32'h001A000F;
14'd558:data <=32'h001C000E;14'd559:data <=32'h001F000F;14'd560:data <=32'h00230011;
14'd561:data <=32'h00290011;14'd562:data <=32'h00320010;14'd563:data <=32'h003C000C;
14'd564:data <=32'h00460003;14'd565:data <=32'h004FFFF7;14'd566:data <=32'h0054FFE8;
14'd567:data <=32'h0056FFD6;14'd568:data <=32'h0052FFC4;14'd569:data <=32'h004BFFB2;
14'd570:data <=32'h0040FFA1;14'd571:data <=32'h0031FF92;14'd572:data <=32'h001EFF85;
14'd573:data <=32'h0007FF7C;14'd574:data <=32'hFFEEFF78;14'd575:data <=32'hFFD2FF7B;
14'd576:data <=32'hFFF8FFD1;14'd577:data <=32'hFFF0FFC6;14'd578:data <=32'hFFE6FFB7;
14'd579:data <=32'hFFBAFF93;14'd580:data <=32'hFF91FFB2;14'd581:data <=32'hFF8BFFCD;
14'd582:data <=32'hFF8BFFE5;14'd583:data <=32'hFF91FFFB;14'd584:data <=32'hFF9B000D;
14'd585:data <=32'hFFA6001A;14'd586:data <=32'hFFB20025;14'd587:data <=32'hFFBF002B;
14'd588:data <=32'hFFCB0030;14'd589:data <=32'hFFD80031;14'd590:data <=32'hFFE3002E;
14'd591:data <=32'hFFEC002A;14'd592:data <=32'hFFF20024;14'd593:data <=32'hFFF4001E;
14'd594:data <=32'hFFF30019;14'd595:data <=32'hFFF10017;14'd596:data <=32'hFFEF0017;
14'd597:data <=32'hFFEE001A;14'd598:data <=32'hFFEF001D;14'd599:data <=32'hFFF2001F;
14'd600:data <=32'hFFF60020;14'd601:data <=32'hFFFA001E;14'd602:data <=32'hFFFD001C;
14'd603:data <=32'hFFFE001A;14'd604:data <=32'hFFFE0017;14'd605:data <=32'hFFFC0017;
14'd606:data <=32'hFFFB0018;14'd607:data <=32'hFFFB001B;14'd608:data <=32'hFFFC001E;
14'd609:data <=32'hFFFE0020;14'd610:data <=32'h00020021;14'd611:data <=32'h00050022;
14'd612:data <=32'h00090022;14'd613:data <=32'h000D0021;14'd614:data <=32'h00100020;
14'd615:data <=32'h0014001F;14'd616:data <=32'h0018001C;14'd617:data <=32'h001B0019;
14'd618:data <=32'h001D0014;14'd619:data <=32'h001E000F;14'd620:data <=32'h001C000A;
14'd621:data <=32'h00170006;14'd622:data <=32'h00120005;14'd623:data <=32'h000B0007;
14'd624:data <=32'h0007000D;14'd625:data <=32'h00060016;14'd626:data <=32'h000A001F;
14'd627:data <=32'h00120028;14'd628:data <=32'h001F002E;14'd629:data <=32'h002E002F;
14'd630:data <=32'h003D002B;14'd631:data <=32'h004D0022;14'd632:data <=32'h00590016;
14'd633:data <=32'h00630005;14'd634:data <=32'h006AFFF2;14'd635:data <=32'h006BFFDD;
14'd636:data <=32'h0069FFC7;14'd637:data <=32'h0060FFB0;14'd638:data <=32'h0052FF9B;
14'd639:data <=32'h003FFF8A;14'd640:data <=32'h0039FFAF;14'd641:data <=32'h002DFF9B;
14'd642:data <=32'h0024FF8E;14'd643:data <=32'h0026FF90;14'd644:data <=32'hFFFAFF99;
14'd645:data <=32'hFFECFFA0;14'd646:data <=32'hFFE1FFA7;14'd647:data <=32'hFFD9FFB0;
14'd648:data <=32'hFFD2FFB7;14'd649:data <=32'hFFCCFFBD;14'd650:data <=32'hFFC5FFC4;
14'd651:data <=32'hFFBEFFCC;14'd652:data <=32'hFFB8FFD6;14'd653:data <=32'hFFB5FFE1;
14'd654:data <=32'hFFB3FFEC;14'd655:data <=32'hFFB3FFF7;14'd656:data <=32'hFFB50001;
14'd657:data <=32'hFFB8000B;14'd658:data <=32'hFFBC0013;14'd659:data <=32'hFFC1001C;
14'd660:data <=32'hFFC70025;14'd661:data <=32'hFFD0002D;14'd662:data <=32'hFFDB0033;
14'd663:data <=32'hFFE80035;14'd664:data <=32'hFFF60034;14'd665:data <=32'h0002002D;
14'd666:data <=32'h000B0023;14'd667:data <=32'h000F0018;14'd668:data <=32'h000E000C;
14'd669:data <=32'h00090002;14'd670:data <=32'h0001FFFC;14'd671:data <=32'hFFF8FFFA;
14'd672:data <=32'hFFF0FFFA;14'd673:data <=32'hFFE9FFFE;14'd674:data <=32'hFFE30004;
14'd675:data <=32'hFFE0000A;14'd676:data <=32'hFFDF0012;14'd677:data <=32'hFFDF001A;
14'd678:data <=32'hFFE10022;14'd679:data <=32'hFFE60029;14'd680:data <=32'hFFED002F;
14'd681:data <=32'hFFF50033;14'd682:data <=32'hFFFF0034;14'd683:data <=32'h00070032;
14'd684:data <=32'h000E002E;14'd685:data <=32'h00120028;14'd686:data <=32'h00130022;
14'd687:data <=32'h0012001E;14'd688:data <=32'h000F001D;14'd689:data <=32'h000D001F;
14'd690:data <=32'h000D0024;14'd691:data <=32'h00100028;14'd692:data <=32'h0015002D;
14'd693:data <=32'h001E002F;14'd694:data <=32'h0028002F;14'd695:data <=32'h0032002C;
14'd696:data <=32'h003B0027;14'd697:data <=32'h0043001F;14'd698:data <=32'h004A0016;
14'd699:data <=32'h004F000C;14'd700:data <=32'h00530001;14'd701:data <=32'h0055FFF4;
14'd702:data <=32'h0054FFE7;14'd703:data <=32'h0050FFD9;14'd704:data <=32'h007BFFF7;
14'd705:data <=32'h0082FFD7;14'd706:data <=32'h0079FFBF;14'd707:data <=32'h0043FFD6;
14'd708:data <=32'h0025FFDB;14'd709:data <=32'h0024FFDD;14'd710:data <=32'h0026FFDC;
14'd711:data <=32'h0029FFD8;14'd712:data <=32'h002BFFD0;14'd713:data <=32'h002AFFC6;
14'd714:data <=32'h0025FFBA;14'd715:data <=32'h001CFFAF;14'd716:data <=32'h000EFFA6;
14'd717:data <=32'hFFFEFFA2;14'd718:data <=32'hFFEDFFA2;14'd719:data <=32'hFFDCFFA5;
14'd720:data <=32'hFFCCFFAC;14'd721:data <=32'hFFBEFFB6;14'd722:data <=32'hFFB1FFC3;
14'd723:data <=32'hFFA8FFD3;14'd724:data <=32'hFFA2FFE6;14'd725:data <=32'hFFA2FFFA;
14'd726:data <=32'hFFA7000F;14'd727:data <=32'hFFB20020;14'd728:data <=32'hFFC2002D;
14'd729:data <=32'hFFD40034;14'd730:data <=32'hFFE60035;14'd731:data <=32'hFFF60030;
14'd732:data <=32'h00020027;14'd733:data <=32'h000A001C;14'd734:data <=32'h000D0010;
14'd735:data <=32'h000C0006;14'd736:data <=32'h0009FFFD;14'd737:data <=32'h0004FFF7;
14'd738:data <=32'hFFFEFFF2;14'd739:data <=32'hFFF7FFEF;14'd740:data <=32'hFFEFFFED;
14'd741:data <=32'hFFE7FFEE;14'd742:data <=32'hFFDFFFF0;14'd743:data <=32'hFFD8FFF6;
14'd744:data <=32'hFFD2FFFD;14'd745:data <=32'hFFCE0006;14'd746:data <=32'hFFCC000F;
14'd747:data <=32'hFFCD0018;14'd748:data <=32'hFFD00020;14'd749:data <=32'hFFD30027;
14'd750:data <=32'hFFD6002E;14'd751:data <=32'hFFD90034;14'd752:data <=32'hFFDD003C;
14'd753:data <=32'hFFE30044;14'd754:data <=32'hFFEC004D;14'd755:data <=32'hFFF80054;
14'd756:data <=32'h00060059;14'd757:data <=32'h00170059;14'd758:data <=32'h00280056;
14'd759:data <=32'h0038004D;14'd760:data <=32'h00440041;14'd761:data <=32'h004C0032;
14'd762:data <=32'h00500023;14'd763:data <=32'h00510015;14'd764:data <=32'h00500008;
14'd765:data <=32'h004BFFFD;14'd766:data <=32'h0046FFF3;14'd767:data <=32'h003FFFEB;
14'd768:data <=32'h00500041;14'd769:data <=32'h00660032;14'd770:data <=32'h00710017;
14'd771:data <=32'h0039FFE7;14'd772:data <=32'h0019FFF1;14'd773:data <=32'h0018FFF9;
14'd774:data <=32'h001C0000;14'd775:data <=32'h00240004;14'd776:data <=32'h002E0004;
14'd777:data <=32'h0038FFFD;14'd778:data <=32'h003FFFF3;14'd779:data <=32'h0043FFE5;
14'd780:data <=32'h0041FFD6;14'd781:data <=32'h003CFFC8;14'd782:data <=32'h0033FFBC;
14'd783:data <=32'h0027FFB2;14'd784:data <=32'h0019FFAB;14'd785:data <=32'h000BFFA7;
14'd786:data <=32'hFFFBFFA6;14'd787:data <=32'hFFEAFFA9;14'd788:data <=32'hFFDAFFAF;
14'd789:data <=32'hFFCCFFBB;14'd790:data <=32'hFFC2FFC9;14'd791:data <=32'hFFBDFFD9;
14'd792:data <=32'hFFBDFFEA;14'd793:data <=32'hFFC1FFF8;14'd794:data <=32'hFFC80003;
14'd795:data <=32'hFFD1000A;14'd796:data <=32'hFFDA000E;14'd797:data <=32'hFFE2000F;
14'd798:data <=32'hFFE80010;14'd799:data <=32'hFFEE000F;14'd800:data <=32'hFFF2000E;
14'd801:data <=32'hFFF7000D;14'd802:data <=32'hFFFD000A;14'd803:data <=32'h00010006;
14'd804:data <=32'h00050000;14'd805:data <=32'h0006FFF9;14'd806:data <=32'h0005FFF0;
14'd807:data <=32'h0001FFE8;14'd808:data <=32'hFFFAFFE2;14'd809:data <=32'hFFF1FFDD;
14'd810:data <=32'hFFE7FFDB;14'd811:data <=32'hFFDCFFDA;14'd812:data <=32'hFFD1FFDD;
14'd813:data <=32'hFFC5FFE2;14'd814:data <=32'hFFBAFFE9;14'd815:data <=32'hFFAFFFF5;
14'd816:data <=32'hFFA60004;14'd817:data <=32'hFFA00017;14'd818:data <=32'hFF9F002D;
14'd819:data <=32'hFFA50043;14'd820:data <=32'hFFB20059;14'd821:data <=32'hFFC4006A;
14'd822:data <=32'hFFDB0076;14'd823:data <=32'hFFF5007B;14'd824:data <=32'h000E0078;
14'd825:data <=32'h00240070;14'd826:data <=32'h00360064;14'd827:data <=32'h00440054;
14'd828:data <=32'h004D0044;14'd829:data <=32'h00520033;14'd830:data <=32'h00540021;
14'd831:data <=32'h00510012;14'd832:data <=32'h00250037;14'd833:data <=32'h00320036;
14'd834:data <=32'h0044002E;14'd835:data <=32'h0057000D;14'd836:data <=32'h0037000B;
14'd837:data <=32'h0033000A;14'd838:data <=32'h00330009;14'd839:data <=32'h0034000A;
14'd840:data <=32'h00380008;14'd841:data <=32'h003D0003;14'd842:data <=32'h0040FFFB;
14'd843:data <=32'h0041FFF2;14'd844:data <=32'h003FFFE8;14'd845:data <=32'h0039FFDE;
14'd846:data <=32'h0033FFD8;14'd847:data <=32'h002BFFD3;14'd848:data <=32'h0024FFD0;
14'd849:data <=32'h001DFFCE;14'd850:data <=32'h0016FFCD;14'd851:data <=32'h0010FFCC;
14'd852:data <=32'h0009FFCC;14'd853:data <=32'h0002FFCF;14'd854:data <=32'hFFFCFFD2;
14'd855:data <=32'hFFF8FFD6;14'd856:data <=32'hFFF6FFDB;14'd857:data <=32'hFFF5FFDF;
14'd858:data <=32'hFFF6FFE1;14'd859:data <=32'hFFF6FFE2;14'd860:data <=32'hFFF5FFE1;
14'd861:data <=32'hFFF2FFE0;14'd862:data <=32'hFFEEFFE1;14'd863:data <=32'hFFE9FFE3;
14'd864:data <=32'hFFE5FFE7;14'd865:data <=32'hFFE2FFEF;14'd866:data <=32'hFFE2FFF6;
14'd867:data <=32'hFFE6FFFD;14'd868:data <=32'hFFEC0002;14'd869:data <=32'hFFF30004;
14'd870:data <=32'hFFFB0003;14'd871:data <=32'h0002FFFF;14'd872:data <=32'h0006FFF9;
14'd873:data <=32'h0009FFF0;14'd874:data <=32'h0008FFE8;14'd875:data <=32'h0006FFDF;
14'd876:data <=32'h0000FFD6;14'd877:data <=32'hFFF7FFCE;14'd878:data <=32'hFFEBFFC7;
14'd879:data <=32'hFFDCFFC4;14'd880:data <=32'hFFCBFFC6;14'd881:data <=32'hFFB9FFCD;
14'd882:data <=32'hFFA9FFD9;14'd883:data <=32'hFF9DFFEB;14'd884:data <=32'hFF960001;
14'd885:data <=32'hFF950017;14'd886:data <=32'hFF9B002D;14'd887:data <=32'hFFA6003F;
14'd888:data <=32'hFFB3004D;14'd889:data <=32'hFFC30057;14'd890:data <=32'hFFD2005D;
14'd891:data <=32'hFFE20060;14'd892:data <=32'hFFF00061;14'd893:data <=32'hFFFD0060;
14'd894:data <=32'h000A005E;14'd895:data <=32'h00170059;14'd896:data <=32'h00240047;
14'd897:data <=32'h002D0042;14'd898:data <=32'h00330041;14'd899:data <=32'h0028005F;
14'd900:data <=32'h001A005F;14'd901:data <=32'h0027005D;14'd902:data <=32'h00350058;
14'd903:data <=32'h00440051;14'd904:data <=32'h00520046;14'd905:data <=32'h005F0037;
14'd906:data <=32'h00680024;14'd907:data <=32'h006A000E;14'd908:data <=32'h0067FFF9;
14'd909:data <=32'h005EFFE5;14'd910:data <=32'h0051FFD6;14'd911:data <=32'h0041FFCD;
14'd912:data <=32'h0031FFC8;14'd913:data <=32'h0022FFC8;14'd914:data <=32'h0015FFCB;
14'd915:data <=32'h000BFFD0;14'd916:data <=32'h0003FFD7;14'd917:data <=32'hFFFDFFDF;
14'd918:data <=32'hFFFAFFE8;14'd919:data <=32'hFFFBFFF0;14'd920:data <=32'hFFFEFFF8;
14'd921:data <=32'h0004FFFE;14'd922:data <=32'h000C0000;14'd923:data <=32'h0014FFFD;
14'd924:data <=32'h001AFFF7;14'd925:data <=32'h001DFFEF;14'd926:data <=32'h001CFFE7;
14'd927:data <=32'h0018FFDF;14'd928:data <=32'h0011FFDB;14'd929:data <=32'h0009FFD9;
14'd930:data <=32'h0002FFDA;14'd931:data <=32'hFFFDFFDD;14'd932:data <=32'hFFFAFFE1;
14'd933:data <=32'hFFF9FFE5;14'd934:data <=32'hFFFAFFE8;14'd935:data <=32'hFFFBFFE9;
14'd936:data <=32'hFFFDFFEA;14'd937:data <=32'hFFFDFFE9;14'd938:data <=32'hFFFEFFE8;
14'd939:data <=32'hFFFFFFE6;14'd940:data <=32'hFFFFFFE2;14'd941:data <=32'hFFFEFFDE;
14'd942:data <=32'hFFFBFFDA;14'd943:data <=32'hFFF7FFD5;14'd944:data <=32'hFFF0FFD1;
14'd945:data <=32'hFFE7FFCF;14'd946:data <=32'hFFDDFFD0;14'd947:data <=32'hFFD3FFD3;
14'd948:data <=32'hFFCBFFD9;14'd949:data <=32'hFFC5FFE1;14'd950:data <=32'hFFC2FFEA;
14'd951:data <=32'hFFC0FFF2;14'd952:data <=32'hFFC0FFF8;14'd953:data <=32'hFFBFFFFC;
14'd954:data <=32'hFFBD0001;14'd955:data <=32'hFFB90006;14'd956:data <=32'hFFB5000E;
14'd957:data <=32'hFFB10018;14'd958:data <=32'hFFB00024;14'd959:data <=32'hFFB10032;
14'd960:data <=32'hFFE4005A;14'd961:data <=32'hFFF0005D;14'd962:data <=32'hFFF50058;
14'd963:data <=32'hFFBE0049;14'd964:data <=32'hFFAE005C;14'd965:data <=32'hFFBD006E;
14'd966:data <=32'hFFD2007D;14'd967:data <=32'hFFEA0087;14'd968:data <=32'h0005008B;
14'd969:data <=32'h00230088;14'd970:data <=32'h003E007C;14'd971:data <=32'h00550069;
14'd972:data <=32'h00650051;14'd973:data <=32'h006E0036;14'd974:data <=32'h006E001C;
14'd975:data <=32'h00680006;14'd976:data <=32'h005EFFF3;14'd977:data <=32'h0051FFE5;
14'd978:data <=32'h0043FFDB;14'd979:data <=32'h0035FFD5;14'd980:data <=32'h0026FFD2;
14'd981:data <=32'h0018FFD4;14'd982:data <=32'h000CFFD8;14'd983:data <=32'h0003FFDF;
14'd984:data <=32'hFFFCFFE9;14'd985:data <=32'hFFFAFFF3;14'd986:data <=32'hFFFCFFFD;
14'd987:data <=32'h00010004;14'd988:data <=32'h00070008;14'd989:data <=32'h000E0009;
14'd990:data <=32'h00130006;14'd991:data <=32'h00170004;14'd992:data <=32'h00190001;
14'd993:data <=32'h001AFFFE;14'd994:data <=32'h001CFFFC;14'd995:data <=32'h001DFFFB;
14'd996:data <=32'h0020FFF8;14'd997:data <=32'h0023FFF5;14'd998:data <=32'h0026FFEF;
14'd999:data <=32'h0027FFE8;14'd1000:data <=32'h0026FFE0;14'd1001:data <=32'h0023FFD8;
14'd1002:data <=32'h001EFFD1;14'd1003:data <=32'h0016FFCB;14'd1004:data <=32'h000EFFC8;
14'd1005:data <=32'h0006FFC6;14'd1006:data <=32'hFFFEFFC6;14'd1007:data <=32'hFFF6FFC7;
14'd1008:data <=32'hFFEEFFC9;14'd1009:data <=32'hFFE7FFCD;14'd1010:data <=32'hFFE1FFD2;
14'd1011:data <=32'hFFDDFFD9;14'd1012:data <=32'hFFDAFFE1;14'd1013:data <=32'hFFDCFFE9;
14'd1014:data <=32'hFFDFFFEE;14'd1015:data <=32'hFFE5FFF1;14'd1016:data <=32'hFFEBFFEF;
14'd1017:data <=32'hFFEEFFEA;14'd1018:data <=32'hFFEEFFE2;14'd1019:data <=32'hFFE9FFDA;
14'd1020:data <=32'hFFE0FFD3;14'd1021:data <=32'hFFD2FFD0;14'd1022:data <=32'hFFC3FFD2;
14'd1023:data <=32'hFFB4FFD9;14'd1024:data <=32'hFFB1000A;14'd1025:data <=32'hFFAD0015;
14'd1026:data <=32'hFFB20018;14'd1027:data <=32'hFFB5FFF6;14'd1028:data <=32'hFF940007;
14'd1029:data <=32'hFF92001B;14'd1030:data <=32'hFF950031;14'd1031:data <=32'hFF9E0046;
14'd1032:data <=32'hFFAD005A;14'd1033:data <=32'hFFC10069;14'd1034:data <=32'hFFD80071;
14'd1035:data <=32'hFFF00073;14'd1036:data <=32'h0006006E;14'd1037:data <=32'h00180065;
14'd1038:data <=32'h00260059;14'd1039:data <=32'h0030004C;14'd1040:data <=32'h00360040;
14'd1041:data <=32'h003A0034;14'd1042:data <=32'h003C0029;14'd1043:data <=32'h003D001F;
14'd1044:data <=32'h003D0014;14'd1045:data <=32'h003A000A;14'd1046:data <=32'h00360001;
14'd1047:data <=32'h0030FFF9;14'd1048:data <=32'h0029FFF5;14'd1049:data <=32'h0022FFF2;
14'd1050:data <=32'h001BFFF1;14'd1051:data <=32'h0016FFF1;14'd1052:data <=32'h0011FFF2;
14'd1053:data <=32'h000DFFF4;14'd1054:data <=32'h0009FFF5;14'd1055:data <=32'h0004FFF8;
14'd1056:data <=32'h0000FFFC;14'd1057:data <=32'hFFFE0002;14'd1058:data <=32'hFFFD000B;
14'd1059:data <=32'h00000013;14'd1060:data <=32'h0008001C;14'd1061:data <=32'h00120021;
14'd1062:data <=32'h001F0022;14'd1063:data <=32'h002C001F;14'd1064:data <=32'h00380017;
14'd1065:data <=32'h0041000B;14'd1066:data <=32'h0046FFFE;14'd1067:data <=32'h0047FFEF;
14'd1068:data <=32'h0045FFE1;14'd1069:data <=32'h003FFFD3;14'd1070:data <=32'h0037FFC8;
14'd1071:data <=32'h002DFFBF;14'd1072:data <=32'h0021FFB9;14'd1073:data <=32'h0013FFB6;
14'd1074:data <=32'h0006FFB5;14'd1075:data <=32'hFFF9FFB9;14'd1076:data <=32'hFFEEFFC0;
14'd1077:data <=32'hFFE7FFC9;14'd1078:data <=32'hFFE4FFD3;14'd1079:data <=32'hFFE5FFDC;
14'd1080:data <=32'hFFEAFFE1;14'd1081:data <=32'hFFEFFFE3;14'd1082:data <=32'hFFF3FFE0;
14'd1083:data <=32'hFFF4FFDA;14'd1084:data <=32'hFFF2FFD3;14'd1085:data <=32'hFFEBFFCD;
14'd1086:data <=32'hFFE1FFCA;14'd1087:data <=32'hFFD7FFC9;14'd1088:data <=32'hFFEEFFC9;
14'd1089:data <=32'hFFDEFFC1;14'd1090:data <=32'hFFD1FFC4;14'd1091:data <=32'hFFD0FFE5;
14'd1092:data <=32'hFFB2FFED;14'd1093:data <=32'hFFAFFFF8;14'd1094:data <=32'hFFAF0004;
14'd1095:data <=32'hFFB1000F;14'd1096:data <=32'hFFB6001B;14'd1097:data <=32'hFFBD0025;
14'd1098:data <=32'hFFC7002C;14'd1099:data <=32'hFFD10030;14'd1100:data <=32'hFFDA0031;
14'd1101:data <=32'hFFE1002F;14'd1102:data <=32'hFFE5002C;14'd1103:data <=32'hFFE6002C;
14'd1104:data <=32'hFFE7002D;14'd1105:data <=32'hFFE80031;14'd1106:data <=32'hFFEB0036;
14'd1107:data <=32'hFFF1003B;14'd1108:data <=32'hFFFA003F;14'd1109:data <=32'h0004003F;
14'd1110:data <=32'h000E003E;14'd1111:data <=32'h0017003A;14'd1112:data <=32'h00200034;
14'd1113:data <=32'h0026002D;14'd1114:data <=32'h002C0025;14'd1115:data <=32'h002F001B;
14'd1116:data <=32'h00300011;14'd1117:data <=32'h002F0006;14'd1118:data <=32'h002AFFFC;
14'd1119:data <=32'h0022FFF3;14'd1120:data <=32'h0017FFEE;14'd1121:data <=32'h000BFFED;
14'd1122:data <=32'hFFFFFFF1;14'd1123:data <=32'hFFF6FFF9;14'd1124:data <=32'hFFF00004;
14'd1125:data <=32'hFFF00011;14'd1126:data <=32'hFFF5001D;14'd1127:data <=32'hFFFD0027;
14'd1128:data <=32'h0009002D;14'd1129:data <=32'h0015002F;14'd1130:data <=32'h0021002D;
14'd1131:data <=32'h002C0029;14'd1132:data <=32'h00350022;14'd1133:data <=32'h003D001A;
14'd1134:data <=32'h00430011;14'd1135:data <=32'h00480006;14'd1136:data <=32'h004AFFFB;
14'd1137:data <=32'h004AFFEF;14'd1138:data <=32'h0047FFE3;14'd1139:data <=32'h0042FFD8;
14'd1140:data <=32'h003BFFD0;14'd1141:data <=32'h0034FFCA;14'd1142:data <=32'h002DFFC5;
14'd1143:data <=32'h0026FFC1;14'd1144:data <=32'h0021FFBE;14'd1145:data <=32'h001CFFB9;
14'd1146:data <=32'h0016FFB3;14'd1147:data <=32'h000EFFAD;14'd1148:data <=32'h0002FFA7;
14'd1149:data <=32'hFFF4FFA4;14'd1150:data <=32'hFFE3FFA5;14'd1151:data <=32'hFFD4FFAA;
14'd1152:data <=32'h001BFFE2;14'd1153:data <=32'h001AFFCF;14'd1154:data <=32'h000BFFBE;
14'd1155:data <=32'hFFC4FFC5;14'd1156:data <=32'hFFA5FFD4;14'd1157:data <=32'hFFA4FFE6;
14'd1158:data <=32'hFFA7FFF7;14'd1159:data <=32'hFFAE0006;14'd1160:data <=32'hFFB70012;
14'd1161:data <=32'hFFC3001B;14'd1162:data <=32'hFFD00020;14'd1163:data <=32'hFFDD0020;
14'd1164:data <=32'hFFE8001B;14'd1165:data <=32'hFFEF0013;14'd1166:data <=32'hFFF1000A;
14'd1167:data <=32'hFFED0002;14'd1168:data <=32'hFFE6FFFD;14'd1169:data <=32'hFFDEFFFD;
14'd1170:data <=32'hFFD60002;14'd1171:data <=32'hFFD0000A;14'd1172:data <=32'hFFCE0014;
14'd1173:data <=32'hFFCF001E;14'd1174:data <=32'hFFD40028;14'd1175:data <=32'hFFDA002F;
14'd1176:data <=32'hFFE30035;14'd1177:data <=32'hFFEB0039;14'd1178:data <=32'hFFF5003B;
14'd1179:data <=32'h0000003C;14'd1180:data <=32'h000B0039;14'd1181:data <=32'h00140033;
14'd1182:data <=32'h001C002A;14'd1183:data <=32'h0020001F;14'd1184:data <=32'h00200015;
14'd1185:data <=32'h001D000B;14'd1186:data <=32'h00170004;14'd1187:data <=32'h000F0001;
14'd1188:data <=32'h00070001;14'd1189:data <=32'h00010004;14'd1190:data <=32'hFFFE0008;
14'd1191:data <=32'hFFFC000D;14'd1192:data <=32'hFFFD0011;14'd1193:data <=32'hFFFE0015;
14'd1194:data <=32'hFFFF0018;14'd1195:data <=32'h0000001B;14'd1196:data <=32'h0001001F;
14'd1197:data <=32'h00040024;14'd1198:data <=32'h00070029;14'd1199:data <=32'h000E002E;
14'd1200:data <=32'h00160032;14'd1201:data <=32'h00200034;14'd1202:data <=32'h002C0034;
14'd1203:data <=32'h00380031;14'd1204:data <=32'h0043002B;14'd1205:data <=32'h004E0023;
14'd1206:data <=32'h00580019;14'd1207:data <=32'h0061000C;14'd1208:data <=32'h006AFFFC;
14'd1209:data <=32'h006FFFE9;14'd1210:data <=32'h0070FFD3;14'd1211:data <=32'h006BFFBB;
14'd1212:data <=32'h0060FFA3;14'd1213:data <=32'h004DFF8F;14'd1214:data <=32'h0035FF80;
14'd1215:data <=32'h0019FF78;14'd1216:data <=32'h001AFFE0;14'd1217:data <=32'h001EFFD3;
14'd1218:data <=32'h0020FFBF;14'd1219:data <=32'h0001FF87;14'd1220:data <=32'hFFD2FF8F;
14'd1221:data <=32'hFFC2FF9F;14'd1222:data <=32'hFFB6FFB1;14'd1223:data <=32'hFFAFFFC3;
14'd1224:data <=32'hFFADFFD7;14'd1225:data <=32'hFFB0FFE8;14'd1226:data <=32'hFFB6FFF8;
14'd1227:data <=32'hFFC10003;14'd1228:data <=32'hFFCD0009;14'd1229:data <=32'hFFD8000B;
14'd1230:data <=32'hFFE00008;14'd1231:data <=32'hFFE50003;14'd1232:data <=32'hFFE5FFFF;
14'd1233:data <=32'hFFE3FFFC;14'd1234:data <=32'hFFDFFFFC;14'd1235:data <=32'hFFDCFFFE;
14'd1236:data <=32'hFFDA0002;14'd1237:data <=32'hFFDA0006;14'd1238:data <=32'hFFDB000A;
14'd1239:data <=32'hFFDD000D;14'd1240:data <=32'hFFDF0010;14'd1241:data <=32'hFFE00012;
14'd1242:data <=32'hFFE20014;14'd1243:data <=32'hFFE40017;14'd1244:data <=32'hFFE6001A;
14'd1245:data <=32'hFFE9001C;14'd1246:data <=32'hFFEE001D;14'd1247:data <=32'hFFF1001D;
14'd1248:data <=32'hFFF3001C;14'd1249:data <=32'hFFF5001B;14'd1250:data <=32'hFFF6001B;
14'd1251:data <=32'hFFF6001B;14'd1252:data <=32'hFFF7001C;14'd1253:data <=32'hFFF9001F;
14'd1254:data <=32'hFFFD0020;14'd1255:data <=32'h00010020;14'd1256:data <=32'h0006001E;
14'd1257:data <=32'h0009001A;14'd1258:data <=32'h000A0014;14'd1259:data <=32'h0008000F;
14'd1260:data <=32'h0004000B;14'd1261:data <=32'hFFFE000A;14'd1262:data <=32'hFFF6000C;
14'd1263:data <=32'hFFF00012;14'd1264:data <=32'hFFED001B;14'd1265:data <=32'hFFEC0025;
14'd1266:data <=32'hFFEF0031;14'd1267:data <=32'hFFF6003C;14'd1268:data <=32'h00000046;
14'd1269:data <=32'h000D004D;14'd1270:data <=32'h001D0053;14'd1271:data <=32'h00300055;
14'd1272:data <=32'h00440052;14'd1273:data <=32'h005A0048;14'd1274:data <=32'h006E0038;
14'd1275:data <=32'h007E0023;14'd1276:data <=32'h00870008;14'd1277:data <=32'h0089FFEB;
14'd1278:data <=32'h0083FFCE;14'd1279:data <=32'h0075FFB5;14'd1280:data <=32'h0053FFDC;
14'd1281:data <=32'h0054FFCA;14'd1282:data <=32'h0058FFBD;14'd1283:data <=32'h0062FFB7;
14'd1284:data <=32'h0039FFAA;14'd1285:data <=32'h002BFFA6;14'd1286:data <=32'h001DFFA3;
14'd1287:data <=32'h0010FFA3;14'd1288:data <=32'h0003FFA5;14'd1289:data <=32'hFFF7FFA9;
14'd1290:data <=32'hFFECFFB0;14'd1291:data <=32'hFFE4FFB7;14'd1292:data <=32'hFFDEFFBD;
14'd1293:data <=32'hFFDAFFC3;14'd1294:data <=32'hFFD6FFC8;14'd1295:data <=32'hFFD0FFCD;
14'd1296:data <=32'hFFCAFFD3;14'd1297:data <=32'hFFC4FFDB;14'd1298:data <=32'hFFBFFFE6;
14'd1299:data <=32'hFFBDFFF3;14'd1300:data <=32'hFFBF0000;14'd1301:data <=32'hFFC6000B;
14'd1302:data <=32'hFFCF0014;14'd1303:data <=32'hFFDA0019;14'd1304:data <=32'hFFE4001A;
14'd1305:data <=32'hFFEE0018;14'd1306:data <=32'hFFF40013;14'd1307:data <=32'hFFF9000D;
14'd1308:data <=32'hFFFB0008;14'd1309:data <=32'hFFFB0002;14'd1310:data <=32'hFFF9FFFD;
14'd1311:data <=32'hFFF6FFF8;14'd1312:data <=32'hFFF1FFF5;14'd1313:data <=32'hFFEBFFF3;
14'd1314:data <=32'hFFE3FFF4;14'd1315:data <=32'hFFDCFFF8;14'd1316:data <=32'hFFD6FFFF;
14'd1317:data <=32'hFFD30008;14'd1318:data <=32'hFFD30012;14'd1319:data <=32'hFFD8001B;
14'd1320:data <=32'hFFDE0021;14'd1321:data <=32'hFFE60025;14'd1322:data <=32'hFFEE0025;
14'd1323:data <=32'hFFF40022;14'd1324:data <=32'hFFF7001D;14'd1325:data <=32'hFFF70019;
14'd1326:data <=32'hFFF50017;14'd1327:data <=32'hFFF20016;14'd1328:data <=32'hFFEE0019;
14'd1329:data <=32'hFFEC001D;14'd1330:data <=32'hFFEA0023;14'd1331:data <=32'hFFEB002A;
14'd1332:data <=32'hFFED0031;14'd1333:data <=32'hFFF10038;14'd1334:data <=32'hFFF70040;
14'd1335:data <=32'h00000047;14'd1336:data <=32'h000C004D;14'd1337:data <=32'h001A0050;
14'd1338:data <=32'h002A004F;14'd1339:data <=32'h003B004A;14'd1340:data <=32'h0049003F;
14'd1341:data <=32'h00550031;14'd1342:data <=32'h005B0021;14'd1343:data <=32'h005E0011;
14'd1344:data <=32'h00700033;14'd1345:data <=32'h0082001E;14'd1346:data <=32'h0086000B;
14'd1347:data <=32'h00560013;14'd1348:data <=32'h003F0009;14'd1349:data <=32'h00440005;
14'd1350:data <=32'h0049FFFE;14'd1351:data <=32'h004DFFF5;14'd1352:data <=32'h0050FFEA;
14'd1353:data <=32'h004FFFDD;14'd1354:data <=32'h004DFFD1;14'd1355:data <=32'h0047FFC5;
14'd1356:data <=32'h0040FFB8;14'd1357:data <=32'h0036FFAC;14'd1358:data <=32'h0028FFA2;
14'd1359:data <=32'h0017FF9A;14'd1360:data <=32'h0003FF96;14'd1361:data <=32'hFFEEFF96;
14'd1362:data <=32'hFFD8FF9E;14'd1363:data <=32'hFFC6FFAC;14'd1364:data <=32'hFFB8FFBE;
14'd1365:data <=32'hFFB1FFD3;14'd1366:data <=32'hFFB1FFE8;14'd1367:data <=32'hFFB7FFFA;
14'd1368:data <=32'hFFC10009;14'd1369:data <=32'hFFCD0013;14'd1370:data <=32'hFFD90019;
14'd1371:data <=32'hFFE6001A;14'd1372:data <=32'hFFF10019;14'd1373:data <=32'hFFFB0015;
14'd1374:data <=32'h0004000F;14'd1375:data <=32'h00090006;14'd1376:data <=32'h000CFFFC;
14'd1377:data <=32'h000BFFF3;14'd1378:data <=32'h0007FFE9;14'd1379:data <=32'hFFFFFFE1;
14'd1380:data <=32'hFFF6FFDD;14'd1381:data <=32'hFFECFFDD;14'd1382:data <=32'hFFE3FFE0;
14'd1383:data <=32'hFFDBFFE4;14'd1384:data <=32'hFFD6FFEA;14'd1385:data <=32'hFFD2FFF0;
14'd1386:data <=32'hFFD1FFF5;14'd1387:data <=32'hFFCFFFFA;14'd1388:data <=32'hFFCCFFFE;
14'd1389:data <=32'hFFC90003;14'd1390:data <=32'hFFC50009;14'd1391:data <=32'hFFC30012;
14'd1392:data <=32'hFFC2001C;14'd1393:data <=32'hFFC40027;14'd1394:data <=32'hFFC90032;
14'd1395:data <=32'hFFD0003C;14'd1396:data <=32'hFFD90044;14'd1397:data <=32'hFFE40049;
14'd1398:data <=32'hFFEF004C;14'd1399:data <=32'hFFFA004E;14'd1400:data <=32'h0006004E;
14'd1401:data <=32'h0011004B;14'd1402:data <=32'h001C0047;14'd1403:data <=32'h00260040;
14'd1404:data <=32'h002E0037;14'd1405:data <=32'h0032002C;14'd1406:data <=32'h00330022;
14'd1407:data <=32'h00300018;14'd1408:data <=32'h00230068;14'd1409:data <=32'h003B0067;
14'd1410:data <=32'h004E0058;14'd1411:data <=32'h002B001E;14'd1412:data <=32'h0011001D;
14'd1413:data <=32'h00140025;14'd1414:data <=32'h001C002B;14'd1415:data <=32'h0028002E;
14'd1416:data <=32'h0033002C;14'd1417:data <=32'h003F0028;14'd1418:data <=32'h004A001F;
14'd1419:data <=32'h00540014;14'd1420:data <=32'h005B0007;14'd1421:data <=32'h0060FFF6;
14'd1422:data <=32'h0060FFE4;14'd1423:data <=32'h005CFFD0;14'd1424:data <=32'h0052FFBD;
14'd1425:data <=32'h0042FFAD;14'd1426:data <=32'h002FFFA3;14'd1427:data <=32'h0019FF9F;
14'd1428:data <=32'h0004FFA1;14'd1429:data <=32'hFFF2FFA9;14'd1430:data <=32'hFFE4FFB4;
14'd1431:data <=32'hFFDAFFC1;14'd1432:data <=32'hFFD5FFCF;14'd1433:data <=32'hFFD3FFDB;
14'd1434:data <=32'hFFD4FFE6;14'd1435:data <=32'hFFD6FFEF;14'd1436:data <=32'hFFD9FFF8;
14'd1437:data <=32'hFFDEFFFF;14'd1438:data <=32'hFFE50006;14'd1439:data <=32'hFFED0009;
14'd1440:data <=32'hFFF5000A;14'd1441:data <=32'hFFFE0009;14'd1442:data <=32'h00050005;
14'd1443:data <=32'h000AFFFF;14'd1444:data <=32'h000DFFF8;14'd1445:data <=32'h000EFFF1;
14'd1446:data <=32'h000DFFEB;14'd1447:data <=32'h000CFFE4;14'd1448:data <=32'h0009FFDE;
14'd1449:data <=32'h0005FFD6;14'd1450:data <=32'h0000FFCF;14'd1451:data <=32'hFFF7FFC8;
14'd1452:data <=32'hFFEBFFC2;14'd1453:data <=32'hFFDCFFBF;14'd1454:data <=32'hFFCBFFC0;
14'd1455:data <=32'hFFBAFFC8;14'd1456:data <=32'hFFA9FFD4;14'd1457:data <=32'hFF9DFFE5;
14'd1458:data <=32'hFF96FFF9;14'd1459:data <=32'hFF94000F;14'd1460:data <=32'hFF980025;
14'd1461:data <=32'hFFA10038;14'd1462:data <=32'hFFAE0049;14'd1463:data <=32'hFFBD0055;
14'd1464:data <=32'hFFCE005E;14'd1465:data <=32'hFFE10063;14'd1466:data <=32'hFFF40064;
14'd1467:data <=32'h00070060;14'd1468:data <=32'h00170056;14'd1469:data <=32'h0023004A;
14'd1470:data <=32'h002A003B;14'd1471:data <=32'h002C002C;14'd1472:data <=32'hFFF4003F;
14'd1473:data <=32'hFFFB0048;14'd1474:data <=32'h000C004C;14'd1475:data <=32'h002A0033;
14'd1476:data <=32'h0010002B;14'd1477:data <=32'h0012002E;14'd1478:data <=32'h00150031;
14'd1479:data <=32'h001B0032;14'd1480:data <=32'h00230032;14'd1481:data <=32'h002A002E;
14'd1482:data <=32'h0030002A;14'd1483:data <=32'h00370025;14'd1484:data <=32'h003C001F;
14'd1485:data <=32'h00410018;14'd1486:data <=32'h0045000F;14'd1487:data <=32'h00480003;
14'd1488:data <=32'h0048FFF8;14'd1489:data <=32'h0044FFEC;14'd1490:data <=32'h003DFFE2;
14'd1491:data <=32'h0034FFDB;14'd1492:data <=32'h002AFFD7;14'd1493:data <=32'h0021FFD6;
14'd1494:data <=32'h001AFFD8;14'd1495:data <=32'h0016FFDA;14'd1496:data <=32'h0013FFDB;
14'd1497:data <=32'h0011FFDB;14'd1498:data <=32'h000EFFDA;14'd1499:data <=32'h000AFFD8;
14'd1500:data <=32'h0005FFD7;14'd1501:data <=32'hFFFFFFD8;14'd1502:data <=32'hFFF8FFDB;
14'd1503:data <=32'hFFF4FFE0;14'd1504:data <=32'hFFF0FFE6;14'd1505:data <=32'hFFF0FFEC;
14'd1506:data <=32'hFFF0FFF2;14'd1507:data <=32'hFFF3FFF8;14'd1508:data <=32'hFFF7FFFC;
14'd1509:data <=32'hFFFCFFFF;14'd1510:data <=32'h00020001;14'd1511:data <=32'h00090001;
14'd1512:data <=32'h0011FFFF;14'd1513:data <=32'h001AFFF9;14'd1514:data <=32'h0020FFEF;
14'd1515:data <=32'h0024FFE3;14'd1516:data <=32'h0023FFD3;14'd1517:data <=32'h001DFFC3;
14'd1518:data <=32'h0011FFB5;14'd1519:data <=32'h0000FFAB;14'd1520:data <=32'hFFECFFA6;
14'd1521:data <=32'hFFD7FFA7;14'd1522:data <=32'hFFC2FFAF;14'd1523:data <=32'hFFB1FFBB;
14'd1524:data <=32'hFFA4FFCA;14'd1525:data <=32'hFF9BFFDC;14'd1526:data <=32'hFF96FFEE;
14'd1527:data <=32'hFF950000;14'd1528:data <=32'hFF970013;14'd1529:data <=32'hFF9D0023;
14'd1530:data <=32'hFFA60033;14'd1531:data <=32'hFFB2003F;14'd1532:data <=32'hFFC00048;
14'd1533:data <=32'hFFCF004C;14'd1534:data <=32'hFFDC004D;14'd1535:data <=32'hFFE7004B;
14'd1536:data <=32'hFFF90038;14'd1537:data <=32'hFFFB0037;14'd1538:data <=32'hFFFA003C;
14'd1539:data <=32'hFFE9005B;14'd1540:data <=32'hFFDA005A;14'd1541:data <=32'hFFE80061;
14'd1542:data <=32'hFFF90066;14'd1543:data <=32'h000B0067;14'd1544:data <=32'h001D0062;
14'd1545:data <=32'h002E0059;14'd1546:data <=32'h003A004C;14'd1547:data <=32'h0043003D;
14'd1548:data <=32'h0048002F;14'd1549:data <=32'h004A0020;14'd1550:data <=32'h00490013;
14'd1551:data <=32'h00460006;14'd1552:data <=32'h003FFFFA;14'd1553:data <=32'h0037FFF1;
14'd1554:data <=32'h002CFFEB;14'd1555:data <=32'h0021FFE9;14'd1556:data <=32'h0016FFEA;
14'd1557:data <=32'h000EFFF0;14'd1558:data <=32'h000AFFF8;14'd1559:data <=32'h000A0000;
14'd1560:data <=32'h000F0007;14'd1561:data <=32'h00150009;14'd1562:data <=32'h001D0008;
14'd1563:data <=32'h00220004;14'd1564:data <=32'h0026FFFE;14'd1565:data <=32'h0027FFF6;
14'd1566:data <=32'h0025FFF0;14'd1567:data <=32'h0021FFEA;14'd1568:data <=32'h001CFFE6;
14'd1569:data <=32'h0018FFE4;14'd1570:data <=32'h0012FFE3;14'd1571:data <=32'h000EFFE4;
14'd1572:data <=32'h0009FFE5;14'd1573:data <=32'h0006FFE8;14'd1574:data <=32'h0004FFEC;
14'd1575:data <=32'h0003FFF0;14'd1576:data <=32'h0006FFF5;14'd1577:data <=32'h000AFFF8;
14'd1578:data <=32'h0011FFF9;14'd1579:data <=32'h0018FFF6;14'd1580:data <=32'h001DFFF0;
14'd1581:data <=32'h0022FFE7;14'd1582:data <=32'h0022FFDD;14'd1583:data <=32'h001EFFD2;
14'd1584:data <=32'h0016FFC9;14'd1585:data <=32'h000EFFC2;14'd1586:data <=32'h0003FFBF;
14'd1587:data <=32'hFFFAFFBE;14'd1588:data <=32'hFFF1FFBE;14'd1589:data <=32'hFFE9FFC0;
14'd1590:data <=32'hFFE1FFC1;14'd1591:data <=32'hFFD9FFC2;14'd1592:data <=32'hFFD1FFC5;
14'd1593:data <=32'hFFC8FFC9;14'd1594:data <=32'hFFBFFFCE;14'd1595:data <=32'hFFB6FFD6;
14'd1596:data <=32'hFFB0FFDF;14'd1597:data <=32'hFFA9FFE9;14'd1598:data <=32'hFFA5FFF3;
14'd1599:data <=32'hFFA1FFFE;14'd1600:data <=32'hFFCA0033;14'd1601:data <=32'hFFCF0035;
14'd1602:data <=32'hFFCD0030;14'd1603:data <=32'hFF970016;14'd1604:data <=32'hFF7E0025;
14'd1605:data <=32'hFF850041;14'd1606:data <=32'hFF93005A;14'd1607:data <=32'hFFA8006F;
14'd1608:data <=32'hFFC2007C;14'd1609:data <=32'hFFDF0082;14'd1610:data <=32'hFFFA0081;
14'd1611:data <=32'h0012007A;14'd1612:data <=32'h0027006E;14'd1613:data <=32'h0037005E;
14'd1614:data <=32'h0043004C;14'd1615:data <=32'h004B0039;14'd1616:data <=32'h004D0026;
14'd1617:data <=32'h004B0013;14'd1618:data <=32'h00430002;14'd1619:data <=32'h0038FFF5;
14'd1620:data <=32'h002AFFEE;14'd1621:data <=32'h001CFFEC;14'd1622:data <=32'h000FFFEF;
14'd1623:data <=32'h0006FFF5;14'd1624:data <=32'h0002FFFD;14'd1625:data <=32'h00020006;
14'd1626:data <=32'h0004000C;14'd1627:data <=32'h00080010;14'd1628:data <=32'h000D0011;
14'd1629:data <=32'h00100011;14'd1630:data <=32'h00130011;14'd1631:data <=32'h00160010;
14'd1632:data <=32'h0018000F;14'd1633:data <=32'h001B000E;14'd1634:data <=32'h001F000D;
14'd1635:data <=32'h0022000A;14'd1636:data <=32'h00250007;14'd1637:data <=32'h00270003;
14'd1638:data <=32'h0027FFFE;14'd1639:data <=32'h0028FFFA;14'd1640:data <=32'h0028FFF6;
14'd1641:data <=32'h0027FFF3;14'd1642:data <=32'h0027FFEF;14'd1643:data <=32'h0027FFEB;
14'd1644:data <=32'h0027FFE5;14'd1645:data <=32'h0024FFE0;14'd1646:data <=32'h0020FFDA;
14'd1647:data <=32'h001AFFD5;14'd1648:data <=32'h0013FFD2;14'd1649:data <=32'h000BFFD3;
14'd1650:data <=32'h0005FFD5;14'd1651:data <=32'h0001FFDB;14'd1652:data <=32'h0001FFDF;
14'd1653:data <=32'h0003FFE3;14'd1654:data <=32'h0008FFE3;14'd1655:data <=32'h000CFFE0;
14'd1656:data <=32'h000FFFDA;14'd1657:data <=32'h0010FFD2;14'd1658:data <=32'h000DFFC8;
14'd1659:data <=32'h0007FFBE;14'd1660:data <=32'hFFFDFFB6;14'd1661:data <=32'hFFF2FFAF;
14'd1662:data <=32'hFFE3FFAA;14'd1663:data <=32'hFFD2FFA8;14'd1664:data <=32'hFFC0FFDF;
14'd1665:data <=32'hFFB8FFE0;14'd1666:data <=32'hFFB7FFDF;14'd1667:data <=32'hFFBCFFBA;
14'd1668:data <=32'hFF91FFBF;14'd1669:data <=32'hFF84FFD6;14'd1670:data <=32'hFF7DFFF1;
14'd1671:data <=32'hFF7D000C;14'd1672:data <=32'hFF850026;14'd1673:data <=32'hFF92003A;
14'd1674:data <=32'hFFA3004A;14'd1675:data <=32'hFFB50056;14'd1676:data <=32'hFFC7005C;
14'd1677:data <=32'hFFD9005F;14'd1678:data <=32'hFFEB005F;14'd1679:data <=32'hFFFB005C;
14'd1680:data <=32'h000A0055;14'd1681:data <=32'h0017004C;14'd1682:data <=32'h00200040;
14'd1683:data <=32'h00250034;14'd1684:data <=32'h00270028;14'd1685:data <=32'h0025001E;
14'd1686:data <=32'h00220017;14'd1687:data <=32'h001E0012;14'd1688:data <=32'h001C000F;
14'd1689:data <=32'h001A000C;14'd1690:data <=32'h00190009;14'd1691:data <=32'h00170005;
14'd1692:data <=32'h00140001;14'd1693:data <=32'h000EFFFE;14'd1694:data <=32'h0008FFFE;
14'd1695:data <=32'h0001FFFF;14'd1696:data <=32'hFFFB0004;14'd1697:data <=32'hFFF7000C;
14'd1698:data <=32'hFFF70014;14'd1699:data <=32'hFFFA001D;14'd1700:data <=32'h00000024;
14'd1701:data <=32'h0008002A;14'd1702:data <=32'h0011002C;14'd1703:data <=32'h001B002C;
14'd1704:data <=32'h0025002B;14'd1705:data <=32'h002F0026;14'd1706:data <=32'h00380020;
14'd1707:data <=32'h00400017;14'd1708:data <=32'h0046000B;14'd1709:data <=32'h0049FFFD;
14'd1710:data <=32'h0047FFEF;14'd1711:data <=32'h0042FFE2;14'd1712:data <=32'h0039FFD7;
14'd1713:data <=32'h002DFFD1;14'd1714:data <=32'h0021FFCE;14'd1715:data <=32'h0016FFD1;
14'd1716:data <=32'h000EFFD7;14'd1717:data <=32'h000BFFDD;14'd1718:data <=32'h000BFFE3;
14'd1719:data <=32'h000FFFE7;14'd1720:data <=32'h0014FFE7;14'd1721:data <=32'h0019FFE4;
14'd1722:data <=32'h001CFFDF;14'd1723:data <=32'h001EFFD8;14'd1724:data <=32'h001DFFCF;
14'd1725:data <=32'h001AFFC5;14'd1726:data <=32'h0015FFBC;14'd1727:data <=32'h000DFFB2;
14'd1728:data <=32'h0018FFBF;14'd1729:data <=32'h000EFFAC;14'd1730:data <=32'h0001FFA4;
14'd1731:data <=32'hFFF7FFBB;14'd1732:data <=32'hFFD0FFB3;14'd1733:data <=32'hFFC4FFBC;
14'd1734:data <=32'hFFBAFFC9;14'd1735:data <=32'hFFB5FFD7;14'd1736:data <=32'hFFB3FFE4;
14'd1737:data <=32'hFFB5FFF0;14'd1738:data <=32'hFFB9FFF8;14'd1739:data <=32'hFFBCFFFF;
14'd1740:data <=32'hFFBE0004;14'd1741:data <=32'hFFBF0009;14'd1742:data <=32'hFFC0000F;
14'd1743:data <=32'hFFC10016;14'd1744:data <=32'hFFC4001D;14'd1745:data <=32'hFFC90024;
14'd1746:data <=32'hFFCE002A;14'd1747:data <=32'hFFD4002F;14'd1748:data <=32'hFFDA0033;
14'd1749:data <=32'hFFE10037;14'd1750:data <=32'hFFE9003B;14'd1751:data <=32'hFFF1003E;
14'd1752:data <=32'hFFFC003F;14'd1753:data <=32'h0008003D;14'd1754:data <=32'h00140038;
14'd1755:data <=32'h001E002F;14'd1756:data <=32'h00240023;14'd1757:data <=32'h00260016;
14'd1758:data <=32'h00230008;14'd1759:data <=32'h001BFFFD;14'd1760:data <=32'h0011FFF7;
14'd1761:data <=32'h0005FFF4;14'd1762:data <=32'hFFFAFFF7;14'd1763:data <=32'hFFF1FFFC;
14'd1764:data <=32'hFFEA0005;14'd1765:data <=32'hFFE7000E;14'd1766:data <=32'hFFE70019;
14'd1767:data <=32'hFFE90023;14'd1768:data <=32'hFFEE002D;14'd1769:data <=32'hFFF70035;
14'd1770:data <=32'h0001003C;14'd1771:data <=32'h000D003F;14'd1772:data <=32'h001B003F;
14'd1773:data <=32'h0029003C;14'd1774:data <=32'h00340034;14'd1775:data <=32'h003D002A;
14'd1776:data <=32'h0043001F;14'd1777:data <=32'h00450013;14'd1778:data <=32'h00440009;
14'd1779:data <=32'h00420002;14'd1780:data <=32'h0040FFFD;14'd1781:data <=32'h003FFFF8;
14'd1782:data <=32'h0040FFF4;14'd1783:data <=32'h0041FFEE;14'd1784:data <=32'h0042FFE6;
14'd1785:data <=32'h0041FFDD;14'd1786:data <=32'h003FFFD3;14'd1787:data <=32'h003AFFC9;
14'd1788:data <=32'h0032FFC1;14'd1789:data <=32'h0029FFB9;14'd1790:data <=32'h0020FFB4;
14'd1791:data <=32'h0015FFB0;14'd1792:data <=32'h003FFFF9;14'd1793:data <=32'h004AFFE1;
14'd1794:data <=32'h0045FFC7;14'd1795:data <=32'h0000FFB3;14'd1796:data <=32'hFFDBFFAF;
14'd1797:data <=32'hFFD0FFBC;14'd1798:data <=32'hFFCAFFCB;14'd1799:data <=32'hFFC9FFDA;
14'd1800:data <=32'hFFCDFFE8;14'd1801:data <=32'hFFD5FFF1;14'd1802:data <=32'hFFDEFFF6;
14'd1803:data <=32'hFFE6FFF5;14'd1804:data <=32'hFFEBFFF1;14'd1805:data <=32'hFFEDFFEB;
14'd1806:data <=32'hFFEAFFE5;14'd1807:data <=32'hFFE5FFE1;14'd1808:data <=32'hFFDEFFE1;
14'd1809:data <=32'hFFD6FFE2;14'd1810:data <=32'hFFCFFFE6;14'd1811:data <=32'hFFC8FFEB;
14'd1812:data <=32'hFFC2FFF3;14'd1813:data <=32'hFFBDFFFC;14'd1814:data <=32'hFFBA0008;
14'd1815:data <=32'hFFBB0016;14'd1816:data <=32'hFFC00023;14'd1817:data <=32'hFFC9002F;
14'd1818:data <=32'hFFD60039;14'd1819:data <=32'hFFE5003D;14'd1820:data <=32'hFFF4003C;
14'd1821:data <=32'h00010036;14'd1822:data <=32'h000B002D;14'd1823:data <=32'h00110023;
14'd1824:data <=32'h00120018;14'd1825:data <=32'h0010000F;14'd1826:data <=32'h000C0009;
14'd1827:data <=32'h00060004;14'd1828:data <=32'h00010001;14'd1829:data <=32'hFFFC0001;
14'd1830:data <=32'hFFF60001;14'd1831:data <=32'hFFF10002;14'd1832:data <=32'hFFEC0006;
14'd1833:data <=32'hFFE7000B;14'd1834:data <=32'hFFE40012;14'd1835:data <=32'hFFE20019;
14'd1836:data <=32'hFFE30022;14'd1837:data <=32'hFFE6002B;14'd1838:data <=32'hFFEB0032;
14'd1839:data <=32'hFFF10039;14'd1840:data <=32'hFFF9003E;14'd1841:data <=32'h00010042;
14'd1842:data <=32'h00090046;14'd1843:data <=32'h0013004A;14'd1844:data <=32'h001F004D;
14'd1845:data <=32'h002D004F;14'd1846:data <=32'h003E004D;14'd1847:data <=32'h00510046;
14'd1848:data <=32'h00620039;14'd1849:data <=32'h00700028;14'd1850:data <=32'h007A0012;
14'd1851:data <=32'h007EFFF9;14'd1852:data <=32'h007BFFE1;14'd1853:data <=32'h0073FFCA;
14'd1854:data <=32'h0065FFB7;14'd1855:data <=32'h0055FFA7;14'd1856:data <=32'h002E000A;
14'd1857:data <=32'h003F0000;14'd1858:data <=32'h004FFFE9;14'd1859:data <=32'h0042FFA1;
14'd1860:data <=32'h0014FF92;14'd1861:data <=32'hFFFEFF98;14'd1862:data <=32'hFFECFFA4;
14'd1863:data <=32'hFFDEFFB3;14'd1864:data <=32'hFFD8FFC4;14'd1865:data <=32'hFFD8FFD4;
14'd1866:data <=32'hFFDDFFE0;14'd1867:data <=32'hFFE3FFE7;14'd1868:data <=32'hFFEAFFEA;
14'd1869:data <=32'hFFEFFFE9;14'd1870:data <=32'hFFF2FFE7;14'd1871:data <=32'hFFF3FFE4;
14'd1872:data <=32'hFFF1FFE2;14'd1873:data <=32'hFFEEFFE0;14'd1874:data <=32'hFFEBFFDF;
14'd1875:data <=32'hFFE7FFDF;14'd1876:data <=32'hFFE2FFE0;14'd1877:data <=32'hFFDDFFE1;
14'd1878:data <=32'hFFD7FFE4;14'd1879:data <=32'hFFD2FFEA;14'd1880:data <=32'hFFCEFFF1;
14'd1881:data <=32'hFFCCFFFA;14'd1882:data <=32'hFFCE0003;14'd1883:data <=32'hFFD2000B;
14'd1884:data <=32'hFFD80010;14'd1885:data <=32'hFFDE0012;14'd1886:data <=32'hFFE30012;
14'd1887:data <=32'hFFE70012;14'd1888:data <=32'hFFE90011;14'd1889:data <=32'hFFE90011;
14'd1890:data <=32'hFFEA0012;14'd1891:data <=32'hFFEB0013;14'd1892:data <=32'hFFEE0015;
14'd1893:data <=32'hFFF20016;14'd1894:data <=32'hFFF60015;14'd1895:data <=32'hFFF90012;
14'd1896:data <=32'hFFFC000E;14'd1897:data <=32'hFFFC000A;14'd1898:data <=32'hFFF90005;
14'd1899:data <=32'hFFF50002;14'd1900:data <=32'hFFEF0000;14'd1901:data <=32'hFFE80001;
14'd1902:data <=32'hFFE20002;14'd1903:data <=32'hFFDB0007;14'd1904:data <=32'hFFD4000D;
14'd1905:data <=32'hFFCF0017;14'd1906:data <=32'hFFCA0023;14'd1907:data <=32'hFFC90032;
14'd1908:data <=32'hFFCC0044;14'd1909:data <=32'hFFD50056;14'd1910:data <=32'hFFE50067;
14'd1911:data <=32'hFFFA0074;14'd1912:data <=32'h0014007A;14'd1913:data <=32'h00300079;
14'd1914:data <=32'h004A0070;14'd1915:data <=32'h00610060;14'd1916:data <=32'h0073004B;
14'd1917:data <=32'h007F0033;14'd1918:data <=32'h0085001A;14'd1919:data <=32'h00860000;
14'd1920:data <=32'h004E0016;14'd1921:data <=32'h005C000C;14'd1922:data <=32'h006B0002;
14'd1923:data <=32'h0081FFF6;14'd1924:data <=32'h0062FFD6;14'd1925:data <=32'h0054FFCA;
14'd1926:data <=32'h0047FFC2;14'd1927:data <=32'h0039FFBE;14'd1928:data <=32'h002DFFBD;
14'd1929:data <=32'h0024FFBE;14'd1930:data <=32'h001EFFC0;14'd1931:data <=32'h0018FFBF;
14'd1932:data <=32'h0013FFBE;14'd1933:data <=32'h000CFFBC;14'd1934:data <=32'h0003FFBA;
14'd1935:data <=32'hFFF9FFBB;14'd1936:data <=32'hFFEEFFBF;14'd1937:data <=32'hFFE5FFC5;
14'd1938:data <=32'hFFDFFFCD;14'd1939:data <=32'hFFDBFFD7;14'd1940:data <=32'hFFD9FFDF;
14'd1941:data <=32'hFFD9FFE7;14'd1942:data <=32'hFFDBFFEE;14'd1943:data <=32'hFFDDFFF3;
14'd1944:data <=32'hFFE0FFF8;14'd1945:data <=32'hFFE5FFFD;14'd1946:data <=32'hFFEAFFFF;
14'd1947:data <=32'hFFF00000;14'd1948:data <=32'hFFF5FFFE;14'd1949:data <=32'hFFFAFFFA;
14'd1950:data <=32'hFFFBFFF3;14'd1951:data <=32'hFFF9FFED;14'd1952:data <=32'hFFF4FFE8;
14'd1953:data <=32'hFFEDFFE5;14'd1954:data <=32'hFFE5FFE6;14'd1955:data <=32'hFFDDFFEA;
14'd1956:data <=32'hFFD8FFF1;14'd1957:data <=32'hFFD6FFF9;14'd1958:data <=32'hFFD70001;
14'd1959:data <=32'hFFDB0007;14'd1960:data <=32'hFFDF000B;14'd1961:data <=32'hFFE4000C;
14'd1962:data <=32'hFFE8000B;14'd1963:data <=32'hFFEA000A;14'd1964:data <=32'hFFEC0008;
14'd1965:data <=32'hFFEC0005;14'd1966:data <=32'hFFEA0002;14'd1967:data <=32'hFFE70000;
14'd1968:data <=32'hFFE2FFFF;14'd1969:data <=32'hFFDBFFFF;14'd1970:data <=32'hFFD30002;
14'd1971:data <=32'hFFCA0009;14'd1972:data <=32'hFFC30014;14'd1973:data <=32'hFFBF0022;
14'd1974:data <=32'hFFC00032;14'd1975:data <=32'hFFC60044;14'd1976:data <=32'hFFD20053;
14'd1977:data <=32'hFFE1005E;14'd1978:data <=32'hFFF40064;14'd1979:data <=32'h00060066;
14'd1980:data <=32'h00180063;14'd1981:data <=32'h0027005D;14'd1982:data <=32'h00340055;
14'd1983:data <=32'h003F004C;14'd1984:data <=32'h00420065;14'd1985:data <=32'h005C005E;
14'd1986:data <=32'h006A0053;14'd1987:data <=32'h0045004E;14'd1988:data <=32'h00380038;
14'd1989:data <=32'h003F0033;14'd1990:data <=32'h0046002D;14'd1991:data <=32'h004C0026;
14'd1992:data <=32'h0053001E;14'd1993:data <=32'h005A0014;14'd1994:data <=32'h00610008;
14'd1995:data <=32'h0066FFF9;14'd1996:data <=32'h0067FFE6;14'd1997:data <=32'h0063FFD2;
14'd1998:data <=32'h005AFFBE;14'd1999:data <=32'h004AFFAD;14'd2000:data <=32'h0036FFA2;
14'd2001:data <=32'h0021FF9D;14'd2002:data <=32'h000BFF9E;14'd2003:data <=32'hFFF8FFA4;
14'd2004:data <=32'hFFE8FFAF;14'd2005:data <=32'hFFDCFFBB;14'd2006:data <=32'hFFD4FFC9;
14'd2007:data <=32'hFFCFFFD8;14'd2008:data <=32'hFFCFFFE7;14'd2009:data <=32'hFFD2FFF5;
14'd2010:data <=32'hFFD90001;14'd2011:data <=32'hFFE3000A;14'd2012:data <=32'hFFEF000F;
14'd2013:data <=32'hFFFC000F;14'd2014:data <=32'h0007000A;14'd2015:data <=32'h00100002;
14'd2016:data <=32'h0013FFF7;14'd2017:data <=32'h0013FFEC;14'd2018:data <=32'h000FFFE4;
14'd2019:data <=32'h0008FFDD;14'd2020:data <=32'h0001FFD9;14'd2021:data <=32'hFFFAFFD8;
14'd2022:data <=32'hFFF4FFD9;14'd2023:data <=32'hFFEFFFDA;14'd2024:data <=32'hFFEBFFDB;
14'd2025:data <=32'hFFE6FFDC;14'd2026:data <=32'hFFE2FFDD;14'd2027:data <=32'hFFDDFFDF;
14'd2028:data <=32'hFFD7FFE2;14'd2029:data <=32'hFFD2FFE6;14'd2030:data <=32'hFFCDFFEA;
14'd2031:data <=32'hFFCAFFF0;14'd2032:data <=32'hFFC7FFF6;14'd2033:data <=32'hFFC5FFFC;
14'd2034:data <=32'hFFC30002;14'd2035:data <=32'hFFC10009;14'd2036:data <=32'hFFC00012;
14'd2037:data <=32'hFFC0001C;14'd2038:data <=32'hFFC30026;14'd2039:data <=32'hFFC80031;
14'd2040:data <=32'hFFD10039;14'd2041:data <=32'hFFDD003F;14'd2042:data <=32'hFFE80041;
14'd2043:data <=32'hFFF2003F;14'd2044:data <=32'hFFFA003B;14'd2045:data <=32'hFFFE0036;
14'd2046:data <=32'hFFFF0032;14'd2047:data <=32'hFFFF0030;14'd2048:data <=32'hFFE10071;
14'd2049:data <=32'hFFF8007F;14'd2050:data <=32'h0010007C;14'd2051:data <=32'h0003003D;
14'd2052:data <=32'hFFEF0033;14'd2053:data <=32'hFFF3003C;14'd2054:data <=32'hFFF90044;
14'd2055:data <=32'h0002004C;14'd2056:data <=32'h000F0053;14'd2057:data <=32'h001F0058;
14'd2058:data <=32'h00320057;14'd2059:data <=32'h00460052;14'd2060:data <=32'h00590045;
14'd2061:data <=32'h00690032;14'd2062:data <=32'h0072001B;14'd2063:data <=32'h00740002;
14'd2064:data <=32'h0070FFEA;14'd2065:data <=32'h0065FFD5;14'd2066:data <=32'h0056FFC5;
14'd2067:data <=32'h0045FFBB;14'd2068:data <=32'h0033FFB4;14'd2069:data <=32'h0022FFB2;
14'd2070:data <=32'h0012FFB3;14'd2071:data <=32'h0003FFB8;14'd2072:data <=32'hFFF6FFBF;
14'd2073:data <=32'hFFEBFFC9;14'd2074:data <=32'hFFE4FFD6;14'd2075:data <=32'hFFE1FFE2;
14'd2076:data <=32'hFFE3FFEF;14'd2077:data <=32'hFFE7FFF9;14'd2078:data <=32'hFFEE0001;
14'd2079:data <=32'hFFF70004;14'd2080:data <=32'hFFFF0006;14'd2081:data <=32'h00060004;
14'd2082:data <=32'h000A0002;14'd2083:data <=32'h000FFFFF;14'd2084:data <=32'h0013FFFC;
14'd2085:data <=32'h0016FFF9;14'd2086:data <=32'h001AFFF4;14'd2087:data <=32'h001EFFEE;
14'd2088:data <=32'h0021FFE5;14'd2089:data <=32'h0021FFDA;14'd2090:data <=32'h001EFFCE;
14'd2091:data <=32'h0017FFC2;14'd2092:data <=32'h000BFFB8;14'd2093:data <=32'hFFFEFFB1;
14'd2094:data <=32'hFFEEFFAE;14'd2095:data <=32'hFFDDFFB0;14'd2096:data <=32'hFFCDFFB4;
14'd2097:data <=32'hFFBFFFBD;14'd2098:data <=32'hFFB2FFC8;14'd2099:data <=32'hFFA7FFD6;
14'd2100:data <=32'hFF9FFFE6;14'd2101:data <=32'hFF9BFFF8;14'd2102:data <=32'hFF9B000B;
14'd2103:data <=32'hFFA2001F;14'd2104:data <=32'hFFAC002F;14'd2105:data <=32'hFFBB003B;
14'd2106:data <=32'hFFCD0042;14'd2107:data <=32'hFFDD0043;14'd2108:data <=32'hFFEC003E;
14'd2109:data <=32'hFFF60035;14'd2110:data <=32'hFFFA002C;14'd2111:data <=32'hFFFB0024;
14'd2112:data <=32'hFFC30028;14'd2113:data <=32'hFFC30038;14'd2114:data <=32'hFFD10046;
14'd2115:data <=32'hFFFA0037;14'd2116:data <=32'hFFE50027;14'd2117:data <=32'hFFE5002B;
14'd2118:data <=32'hFFE50031;14'd2119:data <=32'hFFE80037;14'd2120:data <=32'hFFED003F;
14'd2121:data <=32'hFFF40046;14'd2122:data <=32'hFFFE004D;14'd2123:data <=32'h000C0051;
14'd2124:data <=32'h001B0050;14'd2125:data <=32'h002B004B;14'd2126:data <=32'h00380041;
14'd2127:data <=32'h00410034;14'd2128:data <=32'h00460026;14'd2129:data <=32'h00470019;
14'd2130:data <=32'h0045000D;14'd2131:data <=32'h00420004;14'd2132:data <=32'h003EFFFD;
14'd2133:data <=32'h003AFFF7;14'd2134:data <=32'h0036FFF1;14'd2135:data <=32'h0032FFEB;
14'd2136:data <=32'h002DFFE6;14'd2137:data <=32'h0027FFE2;14'd2138:data <=32'h0020FFDF;
14'd2139:data <=32'h0019FFDE;14'd2140:data <=32'h0012FFDF;14'd2141:data <=32'h000DFFE1;
14'd2142:data <=32'h0009FFE3;14'd2143:data <=32'h0005FFE5;14'd2144:data <=32'h0002FFE8;
14'd2145:data <=32'hFFFFFFEB;14'd2146:data <=32'hFFFBFFF0;14'd2147:data <=32'hFFF9FFF6;
14'd2148:data <=32'hFFFAFFFE;14'd2149:data <=32'hFFFD0006;14'd2150:data <=32'h0004000D;
14'd2151:data <=32'h000F0011;14'd2152:data <=32'h001C0011;14'd2153:data <=32'h0029000C;
14'd2154:data <=32'h00350002;14'd2155:data <=32'h003DFFF3;14'd2156:data <=32'h003FFFE3;
14'd2157:data <=32'h003DFFD1;14'd2158:data <=32'h0036FFC0;14'd2159:data <=32'h002BFFB2;
14'd2160:data <=32'h001DFFA7;14'd2161:data <=32'h000BFF9F;14'd2162:data <=32'hFFF9FF9B;
14'd2163:data <=32'hFFE6FF9B;14'd2164:data <=32'hFFD2FF9F;14'd2165:data <=32'hFFC0FFA9;
14'd2166:data <=32'hFFB0FFB7;14'd2167:data <=32'hFFA5FFC8;14'd2168:data <=32'hFF9EFFDB;
14'd2169:data <=32'hFF9EFFEF;14'd2170:data <=32'hFFA30000;14'd2171:data <=32'hFFAB000D;
14'd2172:data <=32'hFFB40016;14'd2173:data <=32'hFFBD001A;14'd2174:data <=32'hFFC4001D;
14'd2175:data <=32'hFFC8001E;14'd2176:data <=32'hFFDD0014;14'd2177:data <=32'hFFD90014;
14'd2178:data <=32'hFFD3001C;14'd2179:data <=32'hFFBF0038;14'd2180:data <=32'hFFB30031;
14'd2181:data <=32'hFFBB003C;14'd2182:data <=32'hFFC60045;14'd2183:data <=32'hFFD2004C;
14'd2184:data <=32'hFFDE0050;14'd2185:data <=32'hFFEA0053;14'd2186:data <=32'hFFF80054;
14'd2187:data <=32'h00050052;14'd2188:data <=32'h0013004D;14'd2189:data <=32'h001F0044;
14'd2190:data <=32'h00280039;14'd2191:data <=32'h002C002B;14'd2192:data <=32'h002C001E;
14'd2193:data <=32'h00280014;14'd2194:data <=32'h0020000D;14'd2195:data <=32'h0019000A;
14'd2196:data <=32'h0012000C;14'd2197:data <=32'h000F000F;14'd2198:data <=32'h000F0013;
14'd2199:data <=32'h00110017;14'd2200:data <=32'h00150018;14'd2201:data <=32'h001A0018;
14'd2202:data <=32'h001E0017;14'd2203:data <=32'h00220014;14'd2204:data <=32'h0025000F;
14'd2205:data <=32'h0028000B;14'd2206:data <=32'h002A0005;14'd2207:data <=32'h002AFFFE;
14'd2208:data <=32'h0028FFF7;14'd2209:data <=32'h0024FFF1;14'd2210:data <=32'h001DFFEC;
14'd2211:data <=32'h0015FFEA;14'd2212:data <=32'h000CFFEC;14'd2213:data <=32'h0006FFF1;
14'd2214:data <=32'h0002FFF9;14'd2215:data <=32'h00020001;14'd2216:data <=32'h00070009;
14'd2217:data <=32'h000F000F;14'd2218:data <=32'h00180011;14'd2219:data <=32'h0023000E;
14'd2220:data <=32'h002B0009;14'd2221:data <=32'h00320001;14'd2222:data <=32'h0036FFF7;
14'd2223:data <=32'h0038FFED;14'd2224:data <=32'h0038FFE3;14'd2225:data <=32'h0036FFD9;
14'd2226:data <=32'h0033FFCF;14'd2227:data <=32'h002DFFC5;14'd2228:data <=32'h0025FFBC;
14'd2229:data <=32'h001BFFB4;14'd2230:data <=32'h0010FFAF;14'd2231:data <=32'h0004FFAC;
14'd2232:data <=32'hFFF8FFAC;14'd2233:data <=32'hFFEDFFAE;14'd2234:data <=32'hFFE4FFB1;
14'd2235:data <=32'hFFDBFFB4;14'd2236:data <=32'hFFD3FFB6;14'd2237:data <=32'hFFC9FFB8;
14'd2238:data <=32'hFFBEFFBC;14'd2239:data <=32'hFFB1FFC2;14'd2240:data <=32'hFFC90006;
14'd2241:data <=32'hFFC90007;14'd2242:data <=32'hFFC60001;14'd2243:data <=32'hFF97FFDC;
14'd2244:data <=32'hFF7CFFE1;14'd2245:data <=32'hFF79FFFB;14'd2246:data <=32'hFF7C0015;
14'd2247:data <=32'hFF85002D;14'd2248:data <=32'hFF920041;14'd2249:data <=32'hFFA30052;
14'd2250:data <=32'hFFB8005F;14'd2251:data <=32'hFFCE0067;14'd2252:data <=32'hFFE60069;
14'd2253:data <=32'hFFFD0065;14'd2254:data <=32'h0011005B;14'd2255:data <=32'h0020004B;
14'd2256:data <=32'h00290039;14'd2257:data <=32'h002B0027;14'd2258:data <=32'h00270017;
14'd2259:data <=32'h001F000C;14'd2260:data <=32'h00160006;14'd2261:data <=32'h000D0004;
14'd2262:data <=32'h00050006;14'd2263:data <=32'h00000009;14'd2264:data <=32'hFFFE000D;
14'd2265:data <=32'hFFFD0011;14'd2266:data <=32'hFFFD0015;14'd2267:data <=32'hFFFE0019;
14'd2268:data <=32'h0001001D;14'd2269:data <=32'h00040020;14'd2270:data <=32'h00090022;
14'd2271:data <=32'h000F0022;14'd2272:data <=32'h00150020;14'd2273:data <=32'h0019001D;
14'd2274:data <=32'h001D0018;14'd2275:data <=32'h001D0013;14'd2276:data <=32'h001D0010;
14'd2277:data <=32'h001B000D;14'd2278:data <=32'h001A000D;14'd2279:data <=32'h001B000E;
14'd2280:data <=32'h001C000E;14'd2281:data <=32'h0020000E;14'd2282:data <=32'h0023000B;
14'd2283:data <=32'h00270008;14'd2284:data <=32'h00280002;14'd2285:data <=32'h0029FFFD;
14'd2286:data <=32'h0027FFF8;14'd2287:data <=32'h0024FFF5;14'd2288:data <=32'h0021FFF4;
14'd2289:data <=32'h001FFFF5;14'd2290:data <=32'h001FFFF6;14'd2291:data <=32'h0021FFF6;
14'd2292:data <=32'h0023FFF6;14'd2293:data <=32'h0027FFF5;14'd2294:data <=32'h002BFFF1;
14'd2295:data <=32'h002EFFEC;14'd2296:data <=32'h0032FFE6;14'd2297:data <=32'h0035FFDE;
14'd2298:data <=32'h0037FFD3;14'd2299:data <=32'h0038FFC7;14'd2300:data <=32'h0035FFB8;
14'd2301:data <=32'h002EFFA7;14'd2302:data <=32'h0021FF96;14'd2303:data <=32'h000DFF89;
14'd2304:data <=32'hFFE2FFC2;14'd2305:data <=32'hFFD9FFBF;14'd2306:data <=32'hFFD9FFBB;
14'd2307:data <=32'hFFE7FF94;14'd2308:data <=32'hFFBEFF89;14'd2309:data <=32'hFFA8FF98;
14'd2310:data <=32'hFF97FFAC;14'd2311:data <=32'hFF8CFFC2;14'd2312:data <=32'hFF85FFDA;
14'd2313:data <=32'hFF83FFF2;14'd2314:data <=32'hFF870009;14'd2315:data <=32'hFF8F001F;
14'd2316:data <=32'hFF9C0031;14'd2317:data <=32'hFFAD003F;14'd2318:data <=32'hFFC10047;
14'd2319:data <=32'hFFD3004A;14'd2320:data <=32'hFFE40047;14'd2321:data <=32'hFFF20040;
14'd2322:data <=32'hFFFA0039;14'd2323:data <=32'hFFFF0031;14'd2324:data <=32'h0002002B;
14'd2325:data <=32'h00040026;14'd2326:data <=32'h00060022;14'd2327:data <=32'h0008001F;
14'd2328:data <=32'h000A001B;14'd2329:data <=32'h000B0016;14'd2330:data <=32'h000A0011;
14'd2331:data <=32'h0009000C;14'd2332:data <=32'h00050009;14'd2333:data <=32'h00000008;
14'd2334:data <=32'hFFFB0008;14'd2335:data <=32'hFFF8000A;14'd2336:data <=32'hFFF5000D;
14'd2337:data <=32'hFFF30011;14'd2338:data <=32'hFFF20015;14'd2339:data <=32'hFFF2001A;
14'd2340:data <=32'hFFF2001F;14'd2341:data <=32'hFFF40025;14'd2342:data <=32'hFFF8002C;
14'd2343:data <=32'hFFFF0032;14'd2344:data <=32'h00080037;14'd2345:data <=32'h00140039;
14'd2346:data <=32'h00200037;14'd2347:data <=32'h002B0031;14'd2348:data <=32'h00350027;
14'd2349:data <=32'h003A001B;14'd2350:data <=32'h003B000F;14'd2351:data <=32'h00370004;
14'd2352:data <=32'h0032FFFC;14'd2353:data <=32'h002BFFF8;14'd2354:data <=32'h0024FFF6;
14'd2355:data <=32'h001FFFF8;14'd2356:data <=32'h001CFFFA;14'd2357:data <=32'h001BFFFE;
14'd2358:data <=32'h001D0001;14'd2359:data <=32'h00200004;14'd2360:data <=32'h00250006;
14'd2361:data <=32'h002C0006;14'd2362:data <=32'h00350004;14'd2363:data <=32'h003FFFFE;
14'd2364:data <=32'h0048FFF3;14'd2365:data <=32'h004FFFE4;14'd2366:data <=32'h0051FFD1;
14'd2367:data <=32'h004DFFBC;14'd2368:data <=32'h0041FFCC;14'd2369:data <=32'h003FFFB5;
14'd2370:data <=32'h0038FFAA;14'd2371:data <=32'h002CFFB9;14'd2372:data <=32'h000CFFA0;
14'd2373:data <=32'hFFFCFFA2;14'd2374:data <=32'hFFEFFFA6;14'd2375:data <=32'hFFE4FFAC;
14'd2376:data <=32'hFFDAFFB3;14'd2377:data <=32'hFFD2FFB9;14'd2378:data <=32'hFFC9FFC1;
14'd2379:data <=32'hFFC3FFCA;14'd2380:data <=32'hFFBEFFD5;14'd2381:data <=32'hFFBBFFDE;
14'd2382:data <=32'hFFBBFFE8;14'd2383:data <=32'hFFBCFFF0;14'd2384:data <=32'hFFBDFFF8;
14'd2385:data <=32'hFFBEFFFD;14'd2386:data <=32'hFFBE0003;14'd2387:data <=32'hFFBE000B;
14'd2388:data <=32'hFFBF0014;14'd2389:data <=32'hFFC2001E;14'd2390:data <=32'hFFC90029;
14'd2391:data <=32'hFFD30031;14'd2392:data <=32'hFFDF0037;14'd2393:data <=32'hFFED0038;
14'd2394:data <=32'hFFFA0035;14'd2395:data <=32'h0005002E;14'd2396:data <=32'h000D0025;
14'd2397:data <=32'h0010001A;14'd2398:data <=32'h00110010;14'd2399:data <=32'h000E0007;
14'd2400:data <=32'h0009FFFF;14'd2401:data <=32'h0003FFFA;14'd2402:data <=32'hFFFAFFF6;
14'd2403:data <=32'hFFF0FFF5;14'd2404:data <=32'hFFE7FFF8;14'd2405:data <=32'hFFDDFFFF;
14'd2406:data <=32'hFFD60008;14'd2407:data <=32'hFFD20015;14'd2408:data <=32'hFFD30022;
14'd2409:data <=32'hFFD80030;14'd2410:data <=32'hFFE2003B;14'd2411:data <=32'hFFEE0042;
14'd2412:data <=32'hFFFC0045;14'd2413:data <=32'h00080044;14'd2414:data <=32'h00130040;
14'd2415:data <=32'h001B003A;14'd2416:data <=32'h00210034;14'd2417:data <=32'h0024002F;
14'd2418:data <=32'h0027002A;14'd2419:data <=32'h002A0027;14'd2420:data <=32'h002D0024;
14'd2421:data <=32'h00310021;14'd2422:data <=32'h0035001C;14'd2423:data <=32'h00380018;
14'd2424:data <=32'h003B0013;14'd2425:data <=32'h003E000E;14'd2426:data <=32'h00410009;
14'd2427:data <=32'h00450003;14'd2428:data <=32'h0049FFFC;14'd2429:data <=32'h004CFFF2;
14'd2430:data <=32'h004DFFE6;14'd2431:data <=32'h004BFFD8;14'd2432:data <=32'h004F0021;
14'd2433:data <=32'h0064000D;14'd2434:data <=32'h0069FFF4;14'd2435:data <=32'h0030FFCD;
14'd2436:data <=32'h0013FFBA;14'd2437:data <=32'h0008FFC0;14'd2438:data <=32'h0001FFC8;
14'd2439:data <=32'hFFFEFFD0;14'd2440:data <=32'hFFFEFFD6;14'd2441:data <=32'h0000FFDA;
14'd2442:data <=32'h0002FFDA;14'd2443:data <=32'h0003FFD9;14'd2444:data <=32'h0004FFD7;
14'd2445:data <=32'h0003FFD4;14'd2446:data <=32'h0001FFCF;14'd2447:data <=32'hFFFDFFCB;
14'd2448:data <=32'hFFF8FFC6;14'd2449:data <=32'hFFEEFFC2;14'd2450:data <=32'hFFE3FFBF;
14'd2451:data <=32'hFFD5FFC1;14'd2452:data <=32'hFFC7FFC7;14'd2453:data <=32'hFFBAFFD3;
14'd2454:data <=32'hFFB2FFE2;14'd2455:data <=32'hFFAEFFF4;14'd2456:data <=32'hFFB10006;
14'd2457:data <=32'hFFB90015;14'd2458:data <=32'hFFC40021;14'd2459:data <=32'hFFD10028;
14'd2460:data <=32'hFFDE002B;14'd2461:data <=32'hFFEA002A;14'd2462:data <=32'hFFF50027;
14'd2463:data <=32'hFFFD0021;14'd2464:data <=32'h0004001A;14'd2465:data <=32'h00070012;
14'd2466:data <=32'h00090009;14'd2467:data <=32'h00080000;14'd2468:data <=32'h0003FFF8;
14'd2469:data <=32'hFFFCFFF2;14'd2470:data <=32'hFFF3FFEF;14'd2471:data <=32'hFFE9FFEF;
14'd2472:data <=32'hFFE0FFF3;14'd2473:data <=32'hFFD9FFF9;14'd2474:data <=32'hFFD40001;
14'd2475:data <=32'hFFD1000A;14'd2476:data <=32'hFFD10011;14'd2477:data <=32'hFFD10019;
14'd2478:data <=32'hFFD1001F;14'd2479:data <=32'hFFD20027;14'd2480:data <=32'hFFD3002F;
14'd2481:data <=32'hFFD50039;14'd2482:data <=32'hFFDA0044;14'd2483:data <=32'hFFE3004F;
14'd2484:data <=32'hFFEE0059;14'd2485:data <=32'hFFFE0061;14'd2486:data <=32'h00100064;
14'd2487:data <=32'h00220064;14'd2488:data <=32'h0035005F;14'd2489:data <=32'h00460056;
14'd2490:data <=32'h0055004A;14'd2491:data <=32'h0061003B;14'd2492:data <=32'h006B002A;
14'd2493:data <=32'h00710016;14'd2494:data <=32'h00730001;14'd2495:data <=32'h0070FFEB;
14'd2496:data <=32'h00250034;14'd2497:data <=32'h003C0033;14'd2498:data <=32'h00530023;
14'd2499:data <=32'h005EFFD9;14'd2500:data <=32'h003CFFBB;14'd2501:data <=32'h0029FFBB;
14'd2502:data <=32'h0019FFC0;14'd2503:data <=32'h000EFFCA;14'd2504:data <=32'h0009FFD2;
14'd2505:data <=32'h0006FFDA;14'd2506:data <=32'h0007FFE0;14'd2507:data <=32'h0008FFE4;
14'd2508:data <=32'h000BFFE6;14'd2509:data <=32'h000EFFE7;14'd2510:data <=32'h0012FFE6;
14'd2511:data <=32'h0015FFE2;14'd2512:data <=32'h0017FFDC;14'd2513:data <=32'h0016FFD4;
14'd2514:data <=32'h0011FFCC;14'd2515:data <=32'h000AFFC5;14'd2516:data <=32'hFFFEFFC0;
14'd2517:data <=32'hFFF1FFC0;14'd2518:data <=32'hFFE5FFC4;14'd2519:data <=32'hFFDBFFCB;
14'd2520:data <=32'hFFD4FFD5;14'd2521:data <=32'hFFD1FFDF;14'd2522:data <=32'hFFD1FFE9;
14'd2523:data <=32'hFFD2FFF1;14'd2524:data <=32'hFFD5FFF6;14'd2525:data <=32'hFFD8FFFB;
14'd2526:data <=32'hFFDAFFFF;14'd2527:data <=32'hFFDD0003;14'd2528:data <=32'hFFE00006;
14'd2529:data <=32'hFFE40009;14'd2530:data <=32'hFFE9000B;14'd2531:data <=32'hFFED000B;
14'd2532:data <=32'hFFF2000A;14'd2533:data <=32'hFFF60007;14'd2534:data <=32'hFFF80003;
14'd2535:data <=32'hFFF90000;14'd2536:data <=32'hFFF8FFFC;14'd2537:data <=32'hFFF7FFF9;
14'd2538:data <=32'hFFF6FFF5;14'd2539:data <=32'hFFF3FFF2;14'd2540:data <=32'hFFEFFFED;
14'd2541:data <=32'hFFE9FFE9;14'd2542:data <=32'hFFE0FFE6;14'd2543:data <=32'hFFD5FFE5;
14'd2544:data <=32'hFFC7FFE8;14'd2545:data <=32'hFFB9FFF1;14'd2546:data <=32'hFFADFFFF;
14'd2547:data <=32'hFFA40012;14'd2548:data <=32'hFFA10028;14'd2549:data <=32'hFFA5003F;
14'd2550:data <=32'hFFAF0055;14'd2551:data <=32'hFFBF0068;14'd2552:data <=32'hFFD40077;
14'd2553:data <=32'hFFEB0080;14'd2554:data <=32'h00030084;14'd2555:data <=32'h001D0083;
14'd2556:data <=32'h0036007C;14'd2557:data <=32'h004D0070;14'd2558:data <=32'h0061005E;
14'd2559:data <=32'h00710048;14'd2560:data <=32'h002D003F;14'd2561:data <=32'h003D003D;
14'd2562:data <=32'h004F003C;14'd2563:data <=32'h006F0035;14'd2564:data <=32'h005D000E;
14'd2565:data <=32'h00570002;14'd2566:data <=32'h0050FFF9;14'd2567:data <=32'h0049FFF3;
14'd2568:data <=32'h0045FFEE;14'd2569:data <=32'h0041FFE9;14'd2570:data <=32'h003DFFE4;
14'd2571:data <=32'h0039FFDE;14'd2572:data <=32'h0033FFD9;14'd2573:data <=32'h002DFFD5;
14'd2574:data <=32'h0026FFD2;14'd2575:data <=32'h0020FFD1;14'd2576:data <=32'h001AFFD0;
14'd2577:data <=32'h0015FFCE;14'd2578:data <=32'h000FFFCE;14'd2579:data <=32'h0009FFCD;
14'd2580:data <=32'h0001FFCE;14'd2581:data <=32'hFFFAFFD1;14'd2582:data <=32'hFFF4FFD7;
14'd2583:data <=32'hFFF0FFDE;14'd2584:data <=32'hFFEFFFE5;14'd2585:data <=32'hFFF1FFEC;
14'd2586:data <=32'hFFF5FFF0;14'd2587:data <=32'hFFFBFFF1;14'd2588:data <=32'hFFFFFFEF;
14'd2589:data <=32'h0001FFEB;14'd2590:data <=32'h0001FFE6;14'd2591:data <=32'hFFFDFFE2;
14'd2592:data <=32'hFFF9FFE0;14'd2593:data <=32'hFFF3FFDF;14'd2594:data <=32'hFFEEFFE1;
14'd2595:data <=32'hFFEAFFE4;14'd2596:data <=32'hFFE8FFE8;14'd2597:data <=32'hFFE6FFEC;
14'd2598:data <=32'hFFE5FFF0;14'd2599:data <=32'hFFE5FFF4;14'd2600:data <=32'hFFE7FFF8;
14'd2601:data <=32'hFFEAFFFB;14'd2602:data <=32'hFFEDFFFC;14'd2603:data <=32'hFFF2FFFB;
14'd2604:data <=32'hFFF7FFF8;14'd2605:data <=32'hFFFAFFF2;14'd2606:data <=32'hFFF9FFEA;
14'd2607:data <=32'hFFF5FFE1;14'd2608:data <=32'hFFECFFDA;14'd2609:data <=32'hFFDFFFD5;
14'd2610:data <=32'hFFD0FFD5;14'd2611:data <=32'hFFC0FFDB;14'd2612:data <=32'hFFB2FFE6;
14'd2613:data <=32'hFFA8FFF5;14'd2614:data <=32'hFFA20007;14'd2615:data <=32'hFFA10019;
14'd2616:data <=32'hFFA5002C;14'd2617:data <=32'hFFAB003C;14'd2618:data <=32'hFFB5004C;
14'd2619:data <=32'hFFC20059;14'd2620:data <=32'hFFD10063;14'd2621:data <=32'hFFE3006A;
14'd2622:data <=32'hFFF5006E;14'd2623:data <=32'h0008006D;14'd2624:data <=32'h00070075;
14'd2625:data <=32'h001F0078;14'd2626:data <=32'h002D0075;14'd2627:data <=32'h0010006A;
14'd2628:data <=32'h000B0052;14'd2629:data <=32'h00130053;14'd2630:data <=32'h001E0054;
14'd2631:data <=32'h00290055;14'd2632:data <=32'h00380052;14'd2633:data <=32'h0048004B;
14'd2634:data <=32'h00560040;14'd2635:data <=32'h0062002F;14'd2636:data <=32'h0069001C;
14'd2637:data <=32'h006B0008;14'd2638:data <=32'h0068FFF4;14'd2639:data <=32'h0061FFE3;
14'd2640:data <=32'h0057FFD3;14'd2641:data <=32'h004AFFC7;14'd2642:data <=32'h003BFFBD;
14'd2643:data <=32'h002BFFB7;14'd2644:data <=32'h0019FFB5;14'd2645:data <=32'h0008FFB8;
14'd2646:data <=32'hFFF8FFC0;14'd2647:data <=32'hFFECFFCC;14'd2648:data <=32'hFFE5FFDB;
14'd2649:data <=32'hFFE4FFEA;14'd2650:data <=32'hFFE8FFF8;14'd2651:data <=32'hFFF10002;
14'd2652:data <=32'hFFFB0007;14'd2653:data <=32'h00060007;14'd2654:data <=32'h000F0004;
14'd2655:data <=32'h0014FFFE;14'd2656:data <=32'h0018FFF7;14'd2657:data <=32'h0019FFF1;
14'd2658:data <=32'h0018FFEB;14'd2659:data <=32'h0016FFE5;14'd2660:data <=32'h0013FFE0;
14'd2661:data <=32'h0010FFDC;14'd2662:data <=32'h000BFFD9;14'd2663:data <=32'h0006FFD7;
14'd2664:data <=32'h0000FFD5;14'd2665:data <=32'hFFFBFFD5;14'd2666:data <=32'hFFF6FFD7;
14'd2667:data <=32'hFFF3FFD9;14'd2668:data <=32'hFFF1FFDB;14'd2669:data <=32'hFFF0FFDB;
14'd2670:data <=32'hFFEEFFDA;14'd2671:data <=32'hFFEBFFD8;14'd2672:data <=32'hFFE6FFD6;
14'd2673:data <=32'hFFE0FFD5;14'd2674:data <=32'hFFD7FFD6;14'd2675:data <=32'hFFCEFFDA;
14'd2676:data <=32'hFFC6FFE1;14'd2677:data <=32'hFFC0FFEB;14'd2678:data <=32'hFFBDFFF5;
14'd2679:data <=32'hFFBDFFFF;14'd2680:data <=32'hFFC00007;14'd2681:data <=32'hFFC3000E;
14'd2682:data <=32'hFFC60013;14'd2683:data <=32'hFFC90017;14'd2684:data <=32'hFFCA001A;
14'd2685:data <=32'hFFCC001F;14'd2686:data <=32'hFFCE0023;14'd2687:data <=32'hFFD00028;
14'd2688:data <=32'hFFAB0058;14'd2689:data <=32'hFFBB006C;14'd2690:data <=32'hFFCF0070;
14'd2691:data <=32'hFFD10031;14'd2692:data <=32'hFFC10023;14'd2693:data <=32'hFFBF0030;
14'd2694:data <=32'hFFC00041;14'd2695:data <=32'hFFC70053;14'd2696:data <=32'hFFD50064;
14'd2697:data <=32'hFFE90070;14'd2698:data <=32'h00010078;14'd2699:data <=32'h001A0077;
14'd2700:data <=32'h00320070;14'd2701:data <=32'h00460063;14'd2702:data <=32'h00570052;
14'd2703:data <=32'h0062003E;14'd2704:data <=32'h00690029;14'd2705:data <=32'h006B0013;
14'd2706:data <=32'h0068FFFE;14'd2707:data <=32'h0061FFEB;14'd2708:data <=32'h0055FFDA;
14'd2709:data <=32'h0045FFCD;14'd2710:data <=32'h0033FFC5;14'd2711:data <=32'h0020FFC3;
14'd2712:data <=32'h000FFFC7;14'd2713:data <=32'h0002FFCF;14'd2714:data <=32'hFFF9FFDA;
14'd2715:data <=32'hFFF5FFE5;14'd2716:data <=32'hFFF4FFF0;14'd2717:data <=32'hFFF7FFF8;
14'd2718:data <=32'hFFFAFFFD;14'd2719:data <=32'hFFFE0002;14'd2720:data <=32'h00020005;
14'd2721:data <=32'h00060008;14'd2722:data <=32'h000B000A;14'd2723:data <=32'h0011000B;
14'd2724:data <=32'h0018000B;14'd2725:data <=32'h00200008;14'd2726:data <=32'h00270003;
14'd2727:data <=32'h002CFFFC;14'd2728:data <=32'h0031FFF3;14'd2729:data <=32'h0032FFE9;
14'd2730:data <=32'h0031FFDF;14'd2731:data <=32'h002EFFD4;14'd2732:data <=32'h002AFFCA;
14'd2733:data <=32'h0023FFC1;14'd2734:data <=32'h001BFFB8;14'd2735:data <=32'h000FFFB1;
14'd2736:data <=32'h0002FFAB;14'd2737:data <=32'hFFF2FFA8;14'd2738:data <=32'hFFE1FFAA;
14'd2739:data <=32'hFFD0FFB0;14'd2740:data <=32'hFFC1FFBC;14'd2741:data <=32'hFFB6FFCB;
14'd2742:data <=32'hFFB1FFDC;14'd2743:data <=32'hFFB1FFED;14'd2744:data <=32'hFFB7FFFC;
14'd2745:data <=32'hFFBE0006;14'd2746:data <=32'hFFC8000D;14'd2747:data <=32'hFFD1000F;
14'd2748:data <=32'hFFD8000F;14'd2749:data <=32'hFFDD000D;14'd2750:data <=32'hFFE0000A;
14'd2751:data <=32'hFFE00006;14'd2752:data <=32'hFFAEFFFD;14'd2753:data <=32'hFFA8000B;
14'd2754:data <=32'hFFAF001A;14'd2755:data <=32'hFFDB0013;14'd2756:data <=32'hFFC9FFFC;
14'd2757:data <=32'hFFC00002;14'd2758:data <=32'hFFB8000D;14'd2759:data <=32'hFFB3001B;
14'd2760:data <=32'hFFB4002C;14'd2761:data <=32'hFFBA003D;14'd2762:data <=32'hFFC6004C;
14'd2763:data <=32'hFFD50056;14'd2764:data <=32'hFFE6005B;14'd2765:data <=32'hFFF7005D;
14'd2766:data <=32'h0006005A;14'd2767:data <=32'h00140055;14'd2768:data <=32'h0020004F;
14'd2769:data <=32'h002A0047;14'd2770:data <=32'h0033003D;14'd2771:data <=32'h003A0032;
14'd2772:data <=32'h003E0026;14'd2773:data <=32'h003F001A;14'd2774:data <=32'h003D000E;
14'd2775:data <=32'h00390005;14'd2776:data <=32'h0033FFFD;14'd2777:data <=32'h002CFFF8;
14'd2778:data <=32'h0027FFF6;14'd2779:data <=32'h0023FFF4;14'd2780:data <=32'h001FFFF2;
14'd2781:data <=32'h001BFFEF;14'd2782:data <=32'h0017FFED;14'd2783:data <=32'h0011FFEC;
14'd2784:data <=32'h000AFFEC;14'd2785:data <=32'h0002FFEF;14'd2786:data <=32'hFFFCFFF6;
14'd2787:data <=32'hFFF8FFFE;14'd2788:data <=32'hFFF80008;14'd2789:data <=32'hFFFC0013;
14'd2790:data <=32'h0003001B;14'd2791:data <=32'h000E0021;14'd2792:data <=32'h001A0023;
14'd2793:data <=32'h00270021;14'd2794:data <=32'h0034001B;14'd2795:data <=32'h003F0013;
14'd2796:data <=32'h00480007;14'd2797:data <=32'h004FFFF9;14'd2798:data <=32'h0053FFE8;
14'd2799:data <=32'h0052FFD5;14'd2800:data <=32'h004CFFC3;14'd2801:data <=32'h0041FFB1;
14'd2802:data <=32'h0030FFA2;14'd2803:data <=32'h001CFF99;14'd2804:data <=32'h0007FF96;
14'd2805:data <=32'hFFF2FF99;14'd2806:data <=32'hFFE0FFA2;14'd2807:data <=32'hFFD2FFAE;
14'd2808:data <=32'hFFCAFFBB;14'd2809:data <=32'hFFC5FFC9;14'd2810:data <=32'hFFC4FFD4;
14'd2811:data <=32'hFFC5FFDD;14'd2812:data <=32'hFFC6FFE4;14'd2813:data <=32'hFFC8FFEA;
14'd2814:data <=32'hFFC9FFEE;14'd2815:data <=32'hFFCBFFF2;14'd2816:data <=32'hFFE1FFF1;
14'd2817:data <=32'hFFDEFFED;14'd2818:data <=32'hFFD6FFF0;14'd2819:data <=32'hFFBD0003;
14'd2820:data <=32'hFFB1FFF2;14'd2821:data <=32'hFFAEFFFC;14'd2822:data <=32'hFFAD0007;
14'd2823:data <=32'hFFAD0014;14'd2824:data <=32'hFFB10022;14'd2825:data <=32'hFFBA002F;
14'd2826:data <=32'hFFC50039;14'd2827:data <=32'hFFD3003F;14'd2828:data <=32'hFFE20040;
14'd2829:data <=32'hFFEE003D;14'd2830:data <=32'hFFF60037;14'd2831:data <=32'hFFFC0031;
14'd2832:data <=32'hFFFF002B;14'd2833:data <=32'h00000027;14'd2834:data <=32'h00000025;
14'd2835:data <=32'h00000024;14'd2836:data <=32'h00010023;14'd2837:data <=32'h00010023;
14'd2838:data <=32'h00030023;14'd2839:data <=32'h00040024;14'd2840:data <=32'h00050026;
14'd2841:data <=32'h00090028;14'd2842:data <=32'h000E0029;14'd2843:data <=32'h0015002A;
14'd2844:data <=32'h001D0027;14'd2845:data <=32'h00240021;14'd2846:data <=32'h00290019;
14'd2847:data <=32'h002B000F;14'd2848:data <=32'h00290004;14'd2849:data <=32'h0023FFFB;
14'd2850:data <=32'h001AFFF6;14'd2851:data <=32'h0011FFF4;14'd2852:data <=32'h0007FFF7;
14'd2853:data <=32'h0000FFFC;14'd2854:data <=32'hFFFD0004;14'd2855:data <=32'hFFFC000D;
14'd2856:data <=32'hFFFF0015;14'd2857:data <=32'h0004001C;14'd2858:data <=32'h000B0022;
14'd2859:data <=32'h00140026;14'd2860:data <=32'h001E0028;14'd2861:data <=32'h00290027;
14'd2862:data <=32'h00350022;14'd2863:data <=32'h0040001A;14'd2864:data <=32'h00490010;
14'd2865:data <=32'h004F0002;14'd2866:data <=32'h0051FFF3;14'd2867:data <=32'h004FFFE4;
14'd2868:data <=32'h0049FFD6;14'd2869:data <=32'h0041FFCC;14'd2870:data <=32'h0039FFC4;
14'd2871:data <=32'h0030FFBF;14'd2872:data <=32'h0029FFBA;14'd2873:data <=32'h0023FFB6;
14'd2874:data <=32'h001BFFB0;14'd2875:data <=32'h0013FFAA;14'd2876:data <=32'h0009FFA5;
14'd2877:data <=32'hFFFCFFA0;14'd2878:data <=32'hFFEDFF9F;14'd2879:data <=32'hFFDEFFA1;
14'd2880:data <=32'hFFDFFFEF;14'd2881:data <=32'hFFE3FFED;14'd2882:data <=32'hFFE5FFE2;
14'd2883:data <=32'hFFC3FFAE;14'd2884:data <=32'hFFA8FFA2;14'd2885:data <=32'hFF99FFB4;
14'd2886:data <=32'hFF8DFFC9;14'd2887:data <=32'hFF86FFE1;14'd2888:data <=32'hFF86FFFA;
14'd2889:data <=32'hFF8C0014;14'd2890:data <=32'hFF990029;14'd2891:data <=32'hFFAC0039;
14'd2892:data <=32'hFFC00043;14'd2893:data <=32'hFFD50044;14'd2894:data <=32'hFFE80040;
14'd2895:data <=32'hFFF60038;14'd2896:data <=32'hFFFE002E;14'd2897:data <=32'h00030024;
14'd2898:data <=32'h0004001B;14'd2899:data <=32'h00020013;14'd2900:data <=32'hFFFF000D;
14'd2901:data <=32'hFFFB000A;14'd2902:data <=32'hFFF60007;14'd2903:data <=32'hFFF00008;
14'd2904:data <=32'hFFEB000B;14'd2905:data <=32'hFFE70011;14'd2906:data <=32'hFFE50018;
14'd2907:data <=32'hFFE80020;14'd2908:data <=32'hFFEC0027;14'd2909:data <=32'hFFF4002C;
14'd2910:data <=32'hFFFD002D;14'd2911:data <=32'h0006002B;14'd2912:data <=32'h000B0026;
14'd2913:data <=32'h000E0021;14'd2914:data <=32'h000F001C;14'd2915:data <=32'h000F0018;
14'd2916:data <=32'h000D0016;14'd2917:data <=32'h000B0016;14'd2918:data <=32'h000B0016;
14'd2919:data <=32'h000C0017;14'd2920:data <=32'h000D0018;14'd2921:data <=32'h000F0018;
14'd2922:data <=32'h00100017;14'd2923:data <=32'h00110017;14'd2924:data <=32'h00120016;
14'd2925:data <=32'h00130017;14'd2926:data <=32'h00140018;14'd2927:data <=32'h0016001A;
14'd2928:data <=32'h001A001A;14'd2929:data <=32'h001E001A;14'd2930:data <=32'h00210019;
14'd2931:data <=32'h00250018;14'd2932:data <=32'h00280017;14'd2933:data <=32'h002C0016;
14'd2934:data <=32'h00320016;14'd2935:data <=32'h003A0015;14'd2936:data <=32'h00440012;
14'd2937:data <=32'h004F000A;14'd2938:data <=32'h005BFFFE;14'd2939:data <=32'h0063FFED;
14'd2940:data <=32'h0066FFD8;14'd2941:data <=32'h0064FFC1;14'd2942:data <=32'h005AFFAA;
14'd2943:data <=32'h004BFF96;14'd2944:data <=32'h0006FFC7;14'd2945:data <=32'h0005FFC3;
14'd2946:data <=32'h000CFFBD;14'd2947:data <=32'h002BFF94;14'd2948:data <=32'h000AFF74;
14'd2949:data <=32'hFFEFFF75;14'd2950:data <=32'hFFD4FF7C;14'd2951:data <=32'hFFBCFF89;
14'd2952:data <=32'hFFA8FF9D;14'd2953:data <=32'hFF9AFFB4;14'd2954:data <=32'hFF94FFCE;
14'd2955:data <=32'hFF95FFE6;14'd2956:data <=32'hFF9CFFFC;14'd2957:data <=32'hFFA7000C;
14'd2958:data <=32'hFFB40017;14'd2959:data <=32'hFFC1001D;14'd2960:data <=32'hFFCC0020;
14'd2961:data <=32'hFFD50020;14'd2962:data <=32'hFFDD0020;14'd2963:data <=32'hFFE4001F;
14'd2964:data <=32'hFFEA001D;14'd2965:data <=32'hFFF0001B;14'd2966:data <=32'hFFF30017;
14'd2967:data <=32'hFFF60013;14'd2968:data <=32'hFFF6000F;14'd2969:data <=32'hFFF5000B;
14'd2970:data <=32'hFFF3000A;14'd2971:data <=32'hFFF1000A;14'd2972:data <=32'hFFF0000B;
14'd2973:data <=32'hFFF0000C;14'd2974:data <=32'hFFF0000C;14'd2975:data <=32'hFFF0000C;
14'd2976:data <=32'hFFEF000B;14'd2977:data <=32'hFFEC000A;14'd2978:data <=32'hFFE8000B;
14'd2979:data <=32'hFFE5000F;14'd2980:data <=32'hFFE20015;14'd2981:data <=32'hFFE1001D;
14'd2982:data <=32'hFFE30026;14'd2983:data <=32'hFFE9002D;14'd2984:data <=32'hFFF10033;
14'd2985:data <=32'hFFFB0036;14'd2986:data <=32'h00050035;14'd2987:data <=32'h000D0032;
14'd2988:data <=32'h0013002D;14'd2989:data <=32'h00180027;14'd2990:data <=32'h001A0021;
14'd2991:data <=32'h001B001C;14'd2992:data <=32'h001A0017;14'd2993:data <=32'h00180014;
14'd2994:data <=32'h00150011;14'd2995:data <=32'h00110011;14'd2996:data <=32'h000D0013;
14'd2997:data <=32'h000A0018;14'd2998:data <=32'h000A0020;14'd2999:data <=32'h000D0029;
14'd3000:data <=32'h00160032;14'd3001:data <=32'h00230038;14'd3002:data <=32'h0034003A;
14'd3003:data <=32'h00470036;14'd3004:data <=32'h0059002A;14'd3005:data <=32'h00670019;
14'd3006:data <=32'h00710004;14'd3007:data <=32'h0074FFED;14'd3008:data <=32'h0053FFF4;
14'd3009:data <=32'h005CFFE4;14'd3010:data <=32'h0060FFDA;14'd3011:data <=32'h005EFFE2;
14'd3012:data <=32'h004EFFBA;14'd3013:data <=32'h0041FFAE;14'd3014:data <=32'h0032FFA6;
14'd3015:data <=32'h0022FFA0;14'd3016:data <=32'h0011FF9F;14'd3017:data <=32'h0001FFA1;
14'd3018:data <=32'hFFF3FFA8;14'd3019:data <=32'hFFE9FFAF;14'd3020:data <=32'hFFE2FFB8;
14'd3021:data <=32'hFFDDFFBE;14'd3022:data <=32'hFFD9FFC4;14'd3023:data <=32'hFFD4FFC8;
14'd3024:data <=32'hFFCFFFCC;14'd3025:data <=32'hFFC8FFD2;14'd3026:data <=32'hFFC2FFDB;
14'd3027:data <=32'hFFBDFFE5;14'd3028:data <=32'hFFBBFFF2;14'd3029:data <=32'hFFBDFFFE;
14'd3030:data <=32'hFFC20009;14'd3031:data <=32'hFFC80012;14'd3032:data <=32'hFFD10019;
14'd3033:data <=32'hFFDA001D;14'd3034:data <=32'hFFE3001F;14'd3035:data <=32'hFFEC001F;
14'd3036:data <=32'hFFF5001D;14'd3037:data <=32'hFFFD0019;14'd3038:data <=32'h00030012;
14'd3039:data <=32'h00070009;14'd3040:data <=32'h0008FFFE;14'd3041:data <=32'h0004FFF4;
14'd3042:data <=32'hFFFCFFEC;14'd3043:data <=32'hFFF1FFE8;14'd3044:data <=32'hFFE4FFE8;
14'd3045:data <=32'hFFD8FFED;14'd3046:data <=32'hFFCEFFF6;14'd3047:data <=32'hFFC90001;
14'd3048:data <=32'hFFC7000E;14'd3049:data <=32'hFFC9001A;14'd3050:data <=32'hFFCF0024;
14'd3051:data <=32'hFFD6002B;14'd3052:data <=32'hFFDE0031;14'd3053:data <=32'hFFE60035;
14'd3054:data <=32'hFFED0036;14'd3055:data <=32'hFFF40037;14'd3056:data <=32'hFFFB0036;
14'd3057:data <=32'h00010035;14'd3058:data <=32'h00060033;14'd3059:data <=32'h00090030;
14'd3060:data <=32'h000B002D;14'd3061:data <=32'h000C002C;14'd3062:data <=32'h000C002D;
14'd3063:data <=32'h000D0030;14'd3064:data <=32'h00110034;14'd3065:data <=32'h00180039;
14'd3066:data <=32'h0022003B;14'd3067:data <=32'h002E003B;14'd3068:data <=32'h003B0035;
14'd3069:data <=32'h0047002D;14'd3070:data <=32'h004F0020;14'd3071:data <=32'h00540013;
14'd3072:data <=32'h0039004D;14'd3073:data <=32'h00550048;14'd3074:data <=32'h00660038;
14'd3075:data <=32'h00430008;14'd3076:data <=32'h0038FFE9;14'd3077:data <=32'h0033FFE6;
14'd3078:data <=32'h002EFFE5;14'd3079:data <=32'h002BFFE4;14'd3080:data <=32'h0028FFE3;
14'd3081:data <=32'h0025FFE4;14'd3082:data <=32'h0025FFE4;14'd3083:data <=32'h0026FFE3;
14'd3084:data <=32'h0029FFE0;14'd3085:data <=32'h002CFFDA;14'd3086:data <=32'h002DFFD1;
14'd3087:data <=32'h002BFFC5;14'd3088:data <=32'h0023FFB9;14'd3089:data <=32'h0017FFAF;
14'd3090:data <=32'h0006FFA8;14'd3091:data <=32'hFFF5FFA7;14'd3092:data <=32'hFFE3FFAC;
14'd3093:data <=32'hFFD3FFB5;14'd3094:data <=32'hFFC8FFC1;14'd3095:data <=32'hFFC0FFD0;
14'd3096:data <=32'hFFBCFFDF;14'd3097:data <=32'hFFBCFFEE;14'd3098:data <=32'hFFBFFFFC;
14'd3099:data <=32'hFFC50008;14'd3100:data <=32'hFFCE0013;14'd3101:data <=32'hFFD9001A;
14'd3102:data <=32'hFFE6001E;14'd3103:data <=32'hFFF4001D;14'd3104:data <=32'hFFFF0017;
14'd3105:data <=32'h0008000E;14'd3106:data <=32'h000C0003;14'd3107:data <=32'h000CFFF8;
14'd3108:data <=32'h0008FFED;14'd3109:data <=32'h0000FFE6;14'd3110:data <=32'hFFF7FFE2;
14'd3111:data <=32'hFFEEFFE1;14'd3112:data <=32'hFFE6FFE2;14'd3113:data <=32'hFFDFFFE5;
14'd3114:data <=32'hFFD9FFE8;14'd3115:data <=32'hFFD3FFEC;14'd3116:data <=32'hFFCDFFF0;
14'd3117:data <=32'hFFC8FFF6;14'd3118:data <=32'hFFC2FFFD;14'd3119:data <=32'hFFBD0006;
14'd3120:data <=32'hFFBA0011;14'd3121:data <=32'hFFB9001D;14'd3122:data <=32'hFFBC0029;
14'd3123:data <=32'hFFC00035;14'd3124:data <=32'hFFC70040;14'd3125:data <=32'hFFCF004A;
14'd3126:data <=32'hFFD90053;14'd3127:data <=32'hFFE5005B;14'd3128:data <=32'hFFF20063;
14'd3129:data <=32'h00030067;14'd3130:data <=32'h00160068;14'd3131:data <=32'h002A0064;
14'd3132:data <=32'h003C005A;14'd3133:data <=32'h004C004C;14'd3134:data <=32'h00570039;
14'd3135:data <=32'h005B0025;14'd3136:data <=32'hFFFA004C;14'd3137:data <=32'h000E0059;
14'd3138:data <=32'h002A005A;14'd3139:data <=32'h00500019;14'd3140:data <=32'h0042FFF4;
14'd3141:data <=32'h0037FFEF;14'd3142:data <=32'h002DFFED;14'd3143:data <=32'h0025FFEF;
14'd3144:data <=32'h001EFFF1;14'd3145:data <=32'h001AFFF6;14'd3146:data <=32'h0018FFFC;
14'd3147:data <=32'h001B0002;14'd3148:data <=32'h00200006;14'd3149:data <=32'h00290007;
14'd3150:data <=32'h00330003;14'd3151:data <=32'h003BFFFA;14'd3152:data <=32'h0040FFED;
14'd3153:data <=32'h003FFFDF;14'd3154:data <=32'h003AFFD1;14'd3155:data <=32'h0030FFC5;
14'd3156:data <=32'h0024FFBE;14'd3157:data <=32'h0016FFBA;14'd3158:data <=32'h000AFFBA;
14'd3159:data <=32'hFFFEFFBC;14'd3160:data <=32'hFFF4FFC0;14'd3161:data <=32'hFFEBFFC6;
14'd3162:data <=32'hFFE4FFCC;14'd3163:data <=32'hFFDEFFD4;14'd3164:data <=32'hFFDAFFDE;
14'd3165:data <=32'hFFD8FFE7;14'd3166:data <=32'hFFDAFFF1;14'd3167:data <=32'hFFDEFFF9;
14'd3168:data <=32'hFFE4FFFF;14'd3169:data <=32'hFFEB0002;14'd3170:data <=32'hFFF10002;
14'd3171:data <=32'hFFF60001;14'd3172:data <=32'hFFF9FFFF;14'd3173:data <=32'hFFFCFFFC;
14'd3174:data <=32'hFFFEFFFA;14'd3175:data <=32'h0000FFF8;14'd3176:data <=32'h0002FFF5;
14'd3177:data <=32'h0005FFF1;14'd3178:data <=32'h0006FFEB;14'd3179:data <=32'h0006FFE2;
14'd3180:data <=32'h0002FFD9;14'd3181:data <=32'hFFFBFFCF;14'd3182:data <=32'hFFEFFFC8;
14'd3183:data <=32'hFFE0FFC4;14'd3184:data <=32'hFFD0FFC4;14'd3185:data <=32'hFFBFFFC9;
14'd3186:data <=32'hFFAEFFD3;14'd3187:data <=32'hFFA1FFE1;14'd3188:data <=32'hFF96FFF3;
14'd3189:data <=32'hFF900007;14'd3190:data <=32'hFF8D001D;14'd3191:data <=32'hFF900034;
14'd3192:data <=32'hFF98004C;14'd3193:data <=32'hFFA60062;14'd3194:data <=32'hFFBA0074;
14'd3195:data <=32'hFFD40081;14'd3196:data <=32'hFFF00086;14'd3197:data <=32'h000C0084;
14'd3198:data <=32'h00250079;14'd3199:data <=32'h00390069;14'd3200:data <=32'hFFF80042;
14'd3201:data <=32'h0001004B;14'd3202:data <=32'h00100058;14'd3203:data <=32'h00370061;
14'd3204:data <=32'h0039003B;14'd3205:data <=32'h003B0030;14'd3206:data <=32'h003B0028;
14'd3207:data <=32'h003B0020;14'd3208:data <=32'h003A0018;14'd3209:data <=32'h00380012;
14'd3210:data <=32'h0035000D;14'd3211:data <=32'h0033000B;14'd3212:data <=32'h00320009;
14'd3213:data <=32'h00330007;14'd3214:data <=32'h00360003;14'd3215:data <=32'h0038FFFD;
14'd3216:data <=32'h0039FFF5;14'd3217:data <=32'h0037FFED;14'd3218:data <=32'h0032FFE5;
14'd3219:data <=32'h002BFFDF;14'd3220:data <=32'h0022FFDB;14'd3221:data <=32'h001AFFDB;
14'd3222:data <=32'h0014FFDE;14'd3223:data <=32'h0010FFE1;14'd3224:data <=32'h000EFFE4;
14'd3225:data <=32'h000DFFE6;14'd3226:data <=32'h000DFFE6;14'd3227:data <=32'h000DFFE6;
14'd3228:data <=32'h000CFFE5;14'd3229:data <=32'h000AFFE4;14'd3230:data <=32'h0008FFE3;
14'd3231:data <=32'h0007FFE3;14'd3232:data <=32'h0005FFE3;14'd3233:data <=32'h0003FFE2;
14'd3234:data <=32'h0000FFE1;14'd3235:data <=32'hFFFCFFE1;14'd3236:data <=32'hFFF9FFE2;
14'd3237:data <=32'hFFF4FFE5;14'd3238:data <=32'hFFF1FFE9;14'd3239:data <=32'hFFF1FFEF;
14'd3240:data <=32'hFFF3FFF6;14'd3241:data <=32'hFFF9FFFB;14'd3242:data <=32'h0000FFFC;
14'd3243:data <=32'h0009FFFA;14'd3244:data <=32'h0011FFF3;14'd3245:data <=32'h0015FFE9;
14'd3246:data <=32'h0015FFDC;14'd3247:data <=32'h0011FFCF;14'd3248:data <=32'h0008FFC4;
14'd3249:data <=32'hFFFBFFBB;14'd3250:data <=32'hFFECFFB6;14'd3251:data <=32'hFFDBFFB5;
14'd3252:data <=32'hFFCBFFB7;14'd3253:data <=32'hFFBAFFBE;14'd3254:data <=32'hFFAAFFC8;
14'd3255:data <=32'hFF9CFFD7;14'd3256:data <=32'hFF92FFEA;14'd3257:data <=32'hFF8CFFFF;
14'd3258:data <=32'hFF8C0016;14'd3259:data <=32'hFF92002C;14'd3260:data <=32'hFF9D0040;
14'd3261:data <=32'hFFAD004F;14'd3262:data <=32'hFFBF0059;14'd3263:data <=32'hFFD0005E;
14'd3264:data <=32'hFFD1005A;14'd3265:data <=32'hFFDE0064;14'd3266:data <=32'hFFE5006A;
14'd3267:data <=32'hFFCC0063;14'd3268:data <=32'hFFD20050;14'd3269:data <=32'hFFDC0058;
14'd3270:data <=32'hFFE9005F;14'd3271:data <=32'hFFF70064;14'd3272:data <=32'h00070065;
14'd3273:data <=32'h00170063;14'd3274:data <=32'h0026005E;14'd3275:data <=32'h00350056;
14'd3276:data <=32'h0041004C;14'd3277:data <=32'h004C0040;14'd3278:data <=32'h00550031;
14'd3279:data <=32'h005B0020;14'd3280:data <=32'h005D000E;14'd3281:data <=32'h005AFFFA;
14'd3282:data <=32'h0051FFE9;14'd3283:data <=32'h0044FFDB;14'd3284:data <=32'h0032FFD3;
14'd3285:data <=32'h0022FFD1;14'd3286:data <=32'h0012FFD4;14'd3287:data <=32'h0007FFDC;
14'd3288:data <=32'h0000FFE6;14'd3289:data <=32'hFFFDFFF0;14'd3290:data <=32'hFFFEFFF9;
14'd3291:data <=32'h0001FFFF;14'd3292:data <=32'h00050004;14'd3293:data <=32'h000B0007;
14'd3294:data <=32'h00110008;14'd3295:data <=32'h00170007;14'd3296:data <=32'h001C0004;
14'd3297:data <=32'h0021FFFF;14'd3298:data <=32'h0024FFF9;14'd3299:data <=32'h0025FFF1;
14'd3300:data <=32'h0023FFE9;14'd3301:data <=32'h001EFFE4;14'd3302:data <=32'h0018FFE0;
14'd3303:data <=32'h0012FFDF;14'd3304:data <=32'h000DFFE0;14'd3305:data <=32'h000BFFE3;
14'd3306:data <=32'h000AFFE6;14'd3307:data <=32'h000CFFE7;14'd3308:data <=32'h000FFFE6;
14'd3309:data <=32'h0011FFE2;14'd3310:data <=32'h0012FFDC;14'd3311:data <=32'h0010FFD6;
14'd3312:data <=32'h000CFFD0;14'd3313:data <=32'h0005FFCB;14'd3314:data <=32'hFFFEFFC8;
14'd3315:data <=32'hFFF6FFC6;14'd3316:data <=32'hFFEEFFC6;14'd3317:data <=32'hFFE7FFC7;
14'd3318:data <=32'hFFDFFFC9;14'd3319:data <=32'hFFD8FFCB;14'd3320:data <=32'hFFD0FFD0;
14'd3321:data <=32'hFFC9FFD5;14'd3322:data <=32'hFFC3FFDC;14'd3323:data <=32'hFFBFFFE4;
14'd3324:data <=32'hFFBDFFED;14'd3325:data <=32'hFFBDFFF4;14'd3326:data <=32'hFFBDFFF9;
14'd3327:data <=32'hFFBCFFFD;14'd3328:data <=32'hFF92001F;14'd3329:data <=32'hFF950032;
14'd3330:data <=32'hFF9E003B;14'd3331:data <=32'hFFAC0004;14'd3332:data <=32'hFFA0FFF6;
14'd3333:data <=32'hFF980008;14'd3334:data <=32'hFF95001D;14'd3335:data <=32'hFF980034;
14'd3336:data <=32'hFFA1004A;14'd3337:data <=32'hFFAF005C;14'd3338:data <=32'hFFC1006B;
14'd3339:data <=32'hFFD60075;14'd3340:data <=32'hFFEC007B;14'd3341:data <=32'h0005007C;
14'd3342:data <=32'h001D0078;14'd3343:data <=32'h0033006D;14'd3344:data <=32'h0047005D;
14'd3345:data <=32'h00550048;14'd3346:data <=32'h005D0030;14'd3347:data <=32'h005D0018;
14'd3348:data <=32'h00560003;14'd3349:data <=32'h004AFFF3;14'd3350:data <=32'h003BFFE7;
14'd3351:data <=32'h002DFFE2;14'd3352:data <=32'h001FFFE1;14'd3353:data <=32'h0014FFE4;
14'd3354:data <=32'h000BFFE8;14'd3355:data <=32'h0005FFED;14'd3356:data <=32'h0000FFF4;
14'd3357:data <=32'hFFFDFFFA;14'd3358:data <=32'hFFFC0001;14'd3359:data <=32'hFFFC0008;
14'd3360:data <=32'hFFFF000F;14'd3361:data <=32'h00040014;14'd3362:data <=32'h000B0018;
14'd3363:data <=32'h00130019;14'd3364:data <=32'h001A0018;14'd3365:data <=32'h00200015;
14'd3366:data <=32'h00250012;14'd3367:data <=32'h002A000D;14'd3368:data <=32'h002E000A;
14'd3369:data <=32'h00320005;14'd3370:data <=32'h0036FFFF;14'd3371:data <=32'h003BFFF7;
14'd3372:data <=32'h003EFFED;14'd3373:data <=32'h003FFFE2;14'd3374:data <=32'h003CFFD4;
14'd3375:data <=32'h0036FFC7;14'd3376:data <=32'h002BFFBC;14'd3377:data <=32'h001EFFB5;
14'd3378:data <=32'h000FFFB2;14'd3379:data <=32'h0000FFB3;14'd3380:data <=32'hFFF4FFB7;
14'd3381:data <=32'hFFEAFFBE;14'd3382:data <=32'hFFE3FFC7;14'd3383:data <=32'hFFDFFFCF;
14'd3384:data <=32'hFFDDFFD6;14'd3385:data <=32'hFFDCFFDE;14'd3386:data <=32'hFFDEFFE4;
14'd3387:data <=32'hFFE1FFE8;14'd3388:data <=32'hFFE5FFEA;14'd3389:data <=32'hFFEAFFEA;
14'd3390:data <=32'hFFEDFFE6;14'd3391:data <=32'hFFEEFFDF;14'd3392:data <=32'hFFBFFFCC;
14'd3393:data <=32'hFFB3FFD0;14'd3394:data <=32'hFFB0FFDD;14'd3395:data <=32'hFFD9FFDF;
14'd3396:data <=32'hFFCAFFC5;14'd3397:data <=32'hFFBAFFCB;14'd3398:data <=32'hFFACFFD7;
14'd3399:data <=32'hFFA1FFE6;14'd3400:data <=32'hFF9BFFF8;14'd3401:data <=32'hFF9A000B;
14'd3402:data <=32'hFF9D001C;14'd3403:data <=32'hFFA2002D;14'd3404:data <=32'hFFAB003D;
14'd3405:data <=32'hFFB8004B;14'd3406:data <=32'hFFC70056;14'd3407:data <=32'hFFD9005D;
14'd3408:data <=32'hFFEC0060;14'd3409:data <=32'hFFFE005D;14'd3410:data <=32'h000F0055;
14'd3411:data <=32'h001B004A;14'd3412:data <=32'h0023003F;14'd3413:data <=32'h00270033;
14'd3414:data <=32'h00280029;14'd3415:data <=32'h00280021;14'd3416:data <=32'h0027001A;
14'd3417:data <=32'h00270015;14'd3418:data <=32'h0026000E;14'd3419:data <=32'h00250008;
14'd3420:data <=32'h00220002;14'd3421:data <=32'h001DFFFC;14'd3422:data <=32'h0016FFF7;
14'd3423:data <=32'h000EFFF5;14'd3424:data <=32'h0006FFF6;14'd3425:data <=32'hFFFFFFFA;
14'd3426:data <=32'hFFFA0000;14'd3427:data <=32'hFFF60006;14'd3428:data <=32'hFFF5000F;
14'd3429:data <=32'hFFF60017;14'd3430:data <=32'hFFF9001F;14'd3431:data <=32'hFFFE0027;
14'd3432:data <=32'h0006002F;14'd3433:data <=32'h00110034;14'd3434:data <=32'h001E0038;
14'd3435:data <=32'h002E0037;14'd3436:data <=32'h003E0031;14'd3437:data <=32'h004E0026;
14'd3438:data <=32'h00590015;14'd3439:data <=32'h00600002;14'd3440:data <=32'h0061FFED;
14'd3441:data <=32'h005BFFDA;14'd3442:data <=32'h0050FFC9;14'd3443:data <=32'h0043FFBC;
14'd3444:data <=32'h0033FFB4;14'd3445:data <=32'h0024FFB0;14'd3446:data <=32'h0016FFB1;
14'd3447:data <=32'h000AFFB3;14'd3448:data <=32'hFFFFFFB7;14'd3449:data <=32'hFFF7FFBD;
14'd3450:data <=32'hFFF0FFC4;14'd3451:data <=32'hFFECFFCB;14'd3452:data <=32'hFFEBFFD2;
14'd3453:data <=32'hFFECFFD8;14'd3454:data <=32'hFFEFFFDA;14'd3455:data <=32'hFFF3FFD9;
14'd3456:data <=32'h0003FFDD;14'd3457:data <=32'h0003FFD1;14'd3458:data <=32'hFFF9FFCB;
14'd3459:data <=32'hFFDBFFD5;14'd3460:data <=32'hFFD2FFBE;14'd3461:data <=32'hFFC6FFC4;
14'd3462:data <=32'hFFBDFFCE;14'd3463:data <=32'hFFB6FFDB;14'd3464:data <=32'hFFB4FFE9;
14'd3465:data <=32'hFFB5FFF5;14'd3466:data <=32'hFFB80000;14'd3467:data <=32'hFFBC0008;
14'd3468:data <=32'hFFC1000F;14'd3469:data <=32'hFFC60014;14'd3470:data <=32'hFFCB0019;
14'd3471:data <=32'hFFD1001D;14'd3472:data <=32'hFFD70020;14'd3473:data <=32'hFFDD0021;
14'd3474:data <=32'hFFE20021;14'd3475:data <=32'hFFE5001F;14'd3476:data <=32'hFFE6001E;
14'd3477:data <=32'hFFE5001F;14'd3478:data <=32'hFFE50021;14'd3479:data <=32'hFFE60026;
14'd3480:data <=32'hFFE9002C;14'd3481:data <=32'hFFEF0032;14'd3482:data <=32'hFFF80036;
14'd3483:data <=32'h00030036;14'd3484:data <=32'h000D0033;14'd3485:data <=32'h0016002C;
14'd3486:data <=32'h001B0023;14'd3487:data <=32'h001E0019;14'd3488:data <=32'h001C000F;
14'd3489:data <=32'h00180007;14'd3490:data <=32'h00130001;14'd3491:data <=32'h000BFFFE;
14'd3492:data <=32'h0004FFFD;14'd3493:data <=32'hFFFCFFFE;14'd3494:data <=32'hFFF50002;
14'd3495:data <=32'hFFEE0009;14'd3496:data <=32'hFFEA0012;14'd3497:data <=32'hFFE9001E;
14'd3498:data <=32'hFFED002A;14'd3499:data <=32'hFFF40036;14'd3500:data <=32'h0000003F;
14'd3501:data <=32'h000F0044;14'd3502:data <=32'h00200044;14'd3503:data <=32'h002F003F;
14'd3504:data <=32'h003D0036;14'd3505:data <=32'h0046002B;14'd3506:data <=32'h004C001F;
14'd3507:data <=32'h004F0013;14'd3508:data <=32'h00500008;14'd3509:data <=32'h0051FFFE;
14'd3510:data <=32'h0050FFF4;14'd3511:data <=32'h004FFFEA;14'd3512:data <=32'h004DFFE0;
14'd3513:data <=32'h004AFFD6;14'd3514:data <=32'h0044FFCC;14'd3515:data <=32'h003DFFC3;
14'd3516:data <=32'h0035FFBC;14'd3517:data <=32'h002CFFB5;14'd3518:data <=32'h0024FFB0;
14'd3519:data <=32'h001BFFAA;14'd3520:data <=32'h0001FFF3;14'd3521:data <=32'h000DFFEE;
14'd3522:data <=32'h0014FFDE;14'd3523:data <=32'h0000FF9E;14'd3524:data <=32'hFFEBFF85;
14'd3525:data <=32'hFFD4FF8D;14'd3526:data <=32'hFFBFFF9C;14'd3527:data <=32'hFFB0FFAF;
14'd3528:data <=32'hFFA7FFC6;14'd3529:data <=32'hFFA5FFDB;14'd3530:data <=32'hFFA9FFEF;
14'd3531:data <=32'hFFB2FFFE;14'd3532:data <=32'hFFBC0009;14'd3533:data <=32'hFFC70011;
14'd3534:data <=32'hFFD20015;14'd3535:data <=32'hFFDC0016;14'd3536:data <=32'hFFE60015;
14'd3537:data <=32'hFFEE0010;14'd3538:data <=32'hFFF3000A;14'd3539:data <=32'hFFF40002;
14'd3540:data <=32'hFFF2FFFB;14'd3541:data <=32'hFFECFFF6;14'd3542:data <=32'hFFE4FFF4;
14'd3543:data <=32'hFFDBFFF7;14'd3544:data <=32'hFFD4FFFD;14'd3545:data <=32'hFFD00007;
14'd3546:data <=32'hFFD00011;14'd3547:data <=32'hFFD4001B;14'd3548:data <=32'hFFDB0022;
14'd3549:data <=32'hFFE30027;14'd3550:data <=32'hFFEB0028;14'd3551:data <=32'hFFF20027;
14'd3552:data <=32'hFFF80025;14'd3553:data <=32'hFFFC0022;14'd3554:data <=32'hFFFF001E;
14'd3555:data <=32'h0001001B;14'd3556:data <=32'h00020018;14'd3557:data <=32'h00030014;
14'd3558:data <=32'h00010011;14'd3559:data <=32'hFFFF000F;14'd3560:data <=32'hFFFB000E;
14'd3561:data <=32'hFFF7000F;14'd3562:data <=32'hFFF40012;14'd3563:data <=32'hFFF20017;
14'd3564:data <=32'hFFF2001D;14'd3565:data <=32'hFFF40022;14'd3566:data <=32'hFFF80026;
14'd3567:data <=32'hFFFD0029;14'd3568:data <=32'h0000002A;14'd3569:data <=32'h0003002C;
14'd3570:data <=32'h0006002E;14'd3571:data <=32'h00080032;14'd3572:data <=32'h000D0036;
14'd3573:data <=32'h0014003C;14'd3574:data <=32'h001E0041;14'd3575:data <=32'h002C0044;
14'd3576:data <=32'h003C0042;14'd3577:data <=32'h004C003C;14'd3578:data <=32'h005C0031;
14'd3579:data <=32'h00690022;14'd3580:data <=32'h00720010;14'd3581:data <=32'h0079FFFD;
14'd3582:data <=32'h007BFFE7;14'd3583:data <=32'h0079FFD0;14'd3584:data <=32'h0020FFE7;
14'd3585:data <=32'h0028FFE4;14'd3586:data <=32'h0038FFDE;14'd3587:data <=32'h0066FFB7;
14'd3588:data <=32'h0054FF89;14'd3589:data <=32'h0037FF7D;14'd3590:data <=32'h001AFF79;
14'd3591:data <=32'hFFFEFF7D;14'd3592:data <=32'hFFE5FF89;14'd3593:data <=32'hFFD3FF99;
14'd3594:data <=32'hFFC7FFAB;14'd3595:data <=32'hFFC0FFBC;14'd3596:data <=32'hFFBDFFCD;
14'd3597:data <=32'hFFBEFFDB;14'd3598:data <=32'hFFC1FFE8;14'd3599:data <=32'hFFC6FFF3;
14'd3600:data <=32'hFFCDFFFC;14'd3601:data <=32'hFFD50002;14'd3602:data <=32'hFFDE0005;
14'd3603:data <=32'hFFE50005;14'd3604:data <=32'hFFEB0002;14'd3605:data <=32'hFFEEFFFE;
14'd3606:data <=32'hFFEEFFF9;14'd3607:data <=32'hFFECFFF7;14'd3608:data <=32'hFFE8FFF7;
14'd3609:data <=32'hFFE5FFF8;14'd3610:data <=32'hFFE4FFFC;14'd3611:data <=32'hFFE4FFFF;
14'd3612:data <=32'hFFE60001;14'd3613:data <=32'hFFE80001;14'd3614:data <=32'hFFE90000;
14'd3615:data <=32'hFFE8FFFF;14'd3616:data <=32'hFFE6FFFE;14'd3617:data <=32'hFFE3FFFE;
14'd3618:data <=32'hFFDF0001;14'd3619:data <=32'hFFDD0005;14'd3620:data <=32'hFFDB000A;
14'd3621:data <=32'hFFDB0010;14'd3622:data <=32'hFFDD0015;14'd3623:data <=32'hFFE0001A;
14'd3624:data <=32'hFFE3001D;14'd3625:data <=32'hFFE70020;14'd3626:data <=32'hFFEB0022;
14'd3627:data <=32'hFFF00024;14'd3628:data <=32'hFFF50024;14'd3629:data <=32'hFFF90023;
14'd3630:data <=32'hFFFE0020;14'd3631:data <=32'h0000001C;14'd3632:data <=32'h00000016;
14'd3633:data <=32'hFFFD0012;14'd3634:data <=32'hFFF70010;14'd3635:data <=32'hFFEF0011;
14'd3636:data <=32'hFFE70018;14'd3637:data <=32'hFFE20022;14'd3638:data <=32'hFFE10030;
14'd3639:data <=32'hFFE6003F;14'd3640:data <=32'hFFF0004D;14'd3641:data <=32'hFFFF0058;
14'd3642:data <=32'h00120060;14'd3643:data <=32'h00250061;14'd3644:data <=32'h003A005E;
14'd3645:data <=32'h004F0056;14'd3646:data <=32'h00620049;14'd3647:data <=32'h00730038;
14'd3648:data <=32'h00490028;14'd3649:data <=32'h005C0021;14'd3650:data <=32'h0069001B;
14'd3651:data <=32'h00710021;14'd3652:data <=32'h0074FFF0;14'd3653:data <=32'h006CFFDC;
14'd3654:data <=32'h0060FFCC;14'd3655:data <=32'h0051FFC0;14'd3656:data <=32'h0042FFB9;
14'd3657:data <=32'h0035FFB6;14'd3658:data <=32'h002AFFB5;14'd3659:data <=32'h0020FFB4;
14'd3660:data <=32'h0017FFB3;14'd3661:data <=32'h000EFFB2;14'd3662:data <=32'h0004FFB3;
14'd3663:data <=32'hFFF9FFB4;14'd3664:data <=32'hFFF0FFB8;14'd3665:data <=32'hFFE6FFBE;
14'd3666:data <=32'hFFDFFFC6;14'd3667:data <=32'hFFDAFFCD;14'd3668:data <=32'hFFD6FFD5;
14'd3669:data <=32'hFFD4FFDD;14'd3670:data <=32'hFFD1FFE4;14'd3671:data <=32'hFFD1FFEC;
14'd3672:data <=32'hFFD1FFF5;14'd3673:data <=32'hFFD4FFFF;14'd3674:data <=32'hFFD90007;
14'd3675:data <=32'hFFE2000D;14'd3676:data <=32'hFFED0010;14'd3677:data <=32'hFFF8000E;
14'd3678:data <=32'h00000009;14'd3679:data <=32'h0006FFFF;14'd3680:data <=32'h0007FFF5;
14'd3681:data <=32'h0005FFEC;14'd3682:data <=32'hFFFDFFE4;14'd3683:data <=32'hFFF5FFDF;
14'd3684:data <=32'hFFEBFFDE;14'd3685:data <=32'hFFE2FFE0;14'd3686:data <=32'hFFD9FFE4;
14'd3687:data <=32'hFFD3FFEA;14'd3688:data <=32'hFFCDFFF2;14'd3689:data <=32'hFFCAFFFA;
14'd3690:data <=32'hFFC90003;14'd3691:data <=32'hFFCA000C;14'd3692:data <=32'hFFCC0015;
14'd3693:data <=32'hFFD2001C;14'd3694:data <=32'hFFD90021;14'd3695:data <=32'hFFE00023;
14'd3696:data <=32'hFFE70022;14'd3697:data <=32'hFFEB001F;14'd3698:data <=32'hFFEC001B;
14'd3699:data <=32'hFFEA0018;14'd3700:data <=32'hFFE50018;14'd3701:data <=32'hFFE0001C;
14'd3702:data <=32'hFFDD0023;14'd3703:data <=32'hFFDC002D;14'd3704:data <=32'hFFDF0038;
14'd3705:data <=32'hFFE60041;14'd3706:data <=32'hFFF00049;14'd3707:data <=32'hFFFB004F;
14'd3708:data <=32'h00080052;14'd3709:data <=32'h00140052;14'd3710:data <=32'h00210051;
14'd3711:data <=32'h002E004D;14'd3712:data <=32'h0008006E;14'd3713:data <=32'h00260078;
14'd3714:data <=32'h003E0073;14'd3715:data <=32'h0032003F;14'd3716:data <=32'h0039001D;
14'd3717:data <=32'h00380016;14'd3718:data <=32'h00360011;14'd3719:data <=32'h0034000E;
14'd3720:data <=32'h0033000E;14'd3721:data <=32'h0035000E;14'd3722:data <=32'h003A000E;
14'd3723:data <=32'h0041000A;14'd3724:data <=32'h00490002;14'd3725:data <=32'h004FFFF7;
14'd3726:data <=32'h0051FFE9;14'd3727:data <=32'h004FFFD9;14'd3728:data <=32'h0048FFCB;
14'd3729:data <=32'h003EFFBE;14'd3730:data <=32'h0032FFB4;14'd3731:data <=32'h0023FFAD;
14'd3732:data <=32'h0013FFAA;14'd3733:data <=32'h0003FFA9;14'd3734:data <=32'hFFF3FFAC;
14'd3735:data <=32'hFFE4FFB4;14'd3736:data <=32'hFFD6FFBE;14'd3737:data <=32'hFFCCFFCE;
14'd3738:data <=32'hFFC8FFDF;14'd3739:data <=32'hFFC8FFF0;14'd3740:data <=32'hFFCFFFFF;
14'd3741:data <=32'hFFDA000B;14'd3742:data <=32'hFFE70011;14'd3743:data <=32'hFFF50012;
14'd3744:data <=32'h0001000E;14'd3745:data <=32'h00090007;14'd3746:data <=32'h000FFFFF;
14'd3747:data <=32'h0010FFF5;14'd3748:data <=32'h0010FFED;14'd3749:data <=32'h000DFFE5;
14'd3750:data <=32'h0009FFDF;14'd3751:data <=32'h0003FFD9;14'd3752:data <=32'hFFFDFFD5;
14'd3753:data <=32'hFFF5FFD1;14'd3754:data <=32'hFFECFFD0;14'd3755:data <=32'hFFE2FFD0;
14'd3756:data <=32'hFFD9FFD4;14'd3757:data <=32'hFFD1FFD9;14'd3758:data <=32'hFFCAFFDF;
14'd3759:data <=32'hFFC4FFE6;14'd3760:data <=32'hFFC0FFED;14'd3761:data <=32'hFFBDFFF4;
14'd3762:data <=32'hFFB9FFFB;14'd3763:data <=32'hFFB60003;14'd3764:data <=32'hFFB2000D;
14'd3765:data <=32'hFFB0001A;14'd3766:data <=32'hFFB10028;14'd3767:data <=32'hFFB50037;
14'd3768:data <=32'hFFBE0046;14'd3769:data <=32'hFFCC0052;14'd3770:data <=32'hFFDC005A;
14'd3771:data <=32'hFFEE005D;14'd3772:data <=32'hFFFE005B;14'd3773:data <=32'h000C0056;
14'd3774:data <=32'h0018004F;14'd3775:data <=32'h00210046;14'd3776:data <=32'hFFC00048;
14'd3777:data <=32'hFFCD0062;14'd3778:data <=32'hFFE90072;14'd3779:data <=32'h00250040;
14'd3780:data <=32'h0029001B;14'd3781:data <=32'h00240013;14'd3782:data <=32'h001B000F;
14'd3783:data <=32'h0013000F;14'd3784:data <=32'h000D0014;14'd3785:data <=32'h000A001D;
14'd3786:data <=32'h000D0026;14'd3787:data <=32'h0015002E;14'd3788:data <=32'h00200032;
14'd3789:data <=32'h002E0031;14'd3790:data <=32'h003C002B;14'd3791:data <=32'h00470021;
14'd3792:data <=32'h004E0014;14'd3793:data <=32'h00520005;14'd3794:data <=32'h0053FFF7;
14'd3795:data <=32'h0050FFE9;14'd3796:data <=32'h004BFFDB;14'd3797:data <=32'h0042FFCF;
14'd3798:data <=32'h0037FFC4;14'd3799:data <=32'h0029FFBD;14'd3800:data <=32'h001AFFB9;
14'd3801:data <=32'h000AFFBA;14'd3802:data <=32'hFFFCFFBF;14'd3803:data <=32'hFFF1FFC8;
14'd3804:data <=32'hFFEAFFD3;14'd3805:data <=32'hFFE7FFDF;14'd3806:data <=32'hFFE8FFE9;
14'd3807:data <=32'hFFEBFFF0;14'd3808:data <=32'hFFEFFFF6;14'd3809:data <=32'hFFF3FFF9;
14'd3810:data <=32'hFFF7FFFC;14'd3811:data <=32'hFFFAFFFE;14'd3812:data <=32'hFFFEFFFF;
14'd3813:data <=32'h00030000;14'd3814:data <=32'h00090000;14'd3815:data <=32'h000FFFFE;
14'd3816:data <=32'h0016FFF9;14'd3817:data <=32'h001BFFF2;14'd3818:data <=32'h001EFFE8;
14'd3819:data <=32'h001EFFDD;14'd3820:data <=32'h001BFFD2;14'd3821:data <=32'h0015FFC7;
14'd3822:data <=32'h000CFFBE;14'd3823:data <=32'h0001FFB6;14'd3824:data <=32'hFFF4FFB0;
14'd3825:data <=32'hFFE4FFAC;14'd3826:data <=32'hFFD2FFAB;14'd3827:data <=32'hFFBFFFAF;
14'd3828:data <=32'hFFACFFB7;14'd3829:data <=32'hFF99FFC6;14'd3830:data <=32'hFF8BFFDA;
14'd3831:data <=32'hFF82FFF3;14'd3832:data <=32'hFF7F000E;14'd3833:data <=32'hFF850029;
14'd3834:data <=32'hFF910040;14'd3835:data <=32'hFFA30053;14'd3836:data <=32'hFFB8005F;
14'd3837:data <=32'hFFCE0066;14'd3838:data <=32'hFFE30067;14'd3839:data <=32'hFFF60063;
14'd3840:data <=32'hFFC80025;14'd3841:data <=32'hFFC70036;14'd3842:data <=32'hFFCF004D;
14'd3843:data <=32'hFFF90066;14'd3844:data <=32'h000B0045;14'd3845:data <=32'h0010003C;
14'd3846:data <=32'h00120033;14'd3847:data <=32'h0011002D;14'd3848:data <=32'h000F002A;
14'd3849:data <=32'h000D002B;14'd3850:data <=32'h000D002D;14'd3851:data <=32'h00110031;
14'd3852:data <=32'h00170032;14'd3853:data <=32'h001F0032;14'd3854:data <=32'h0027002E;
14'd3855:data <=32'h002E0028;14'd3856:data <=32'h00330020;14'd3857:data <=32'h00350018;
14'd3858:data <=32'h00350010;14'd3859:data <=32'h0034000A;14'd3860:data <=32'h00330004;
14'd3861:data <=32'h0031FFFE;14'd3862:data <=32'h0030FFF9;14'd3863:data <=32'h002DFFF4;
14'd3864:data <=32'h0029FFF0;14'd3865:data <=32'h0024FFEC;14'd3866:data <=32'h001FFFEB;
14'd3867:data <=32'h001BFFEB;14'd3868:data <=32'h0018FFEC;14'd3869:data <=32'h0017FFED;
14'd3870:data <=32'h0016FFED;14'd3871:data <=32'h0016FFEB;14'd3872:data <=32'h0015FFE8;
14'd3873:data <=32'h0012FFE5;14'd3874:data <=32'h000DFFE3;14'd3875:data <=32'h0007FFE3;
14'd3876:data <=32'h0001FFE5;14'd3877:data <=32'hFFFCFFEB;14'd3878:data <=32'hFFFAFFF2;
14'd3879:data <=32'hFFFCFFFA;14'd3880:data <=32'h00010001;14'd3881:data <=32'h00080005;
14'd3882:data <=32'h00120006;14'd3883:data <=32'h001B0003;14'd3884:data <=32'h0024FFFD;
14'd3885:data <=32'h002BFFF4;14'd3886:data <=32'h0030FFE9;14'd3887:data <=32'h0031FFDC;
14'd3888:data <=32'h0030FFCD;14'd3889:data <=32'h002BFFBE;14'd3890:data <=32'h0021FFAF;
14'd3891:data <=32'h0012FFA1;14'd3892:data <=32'hFFFFFF98;14'd3893:data <=32'hFFE8FF94;
14'd3894:data <=32'hFFD0FF96;14'd3895:data <=32'hFFB9FF9F;14'd3896:data <=32'hFFA6FFAF;
14'd3897:data <=32'hFF98FFC3;14'd3898:data <=32'hFF90FFD8;14'd3899:data <=32'hFF8EFFEE;
14'd3900:data <=32'hFF910001;14'd3901:data <=32'hFF960012;14'd3902:data <=32'hFF9E0021;
14'd3903:data <=32'hFFA6002C;14'd3904:data <=32'hFFB10026;14'd3905:data <=32'hFFB30034;
14'd3906:data <=32'hFFB3003F;14'd3907:data <=32'hFF9E003A;14'd3908:data <=32'hFFAE002C;
14'd3909:data <=32'hFFB50036;14'd3910:data <=32'hFFBC003F;14'd3911:data <=32'hFFC50048;
14'd3912:data <=32'hFFCE004F;14'd3913:data <=32'hFFD80057;14'd3914:data <=32'hFFE5005E;
14'd3915:data <=32'hFFF50062;14'd3916:data <=32'h00070063;14'd3917:data <=32'h001A005E;
14'd3918:data <=32'h002B0054;14'd3919:data <=32'h00380046;14'd3920:data <=32'h00400035;
14'd3921:data <=32'h00420024;14'd3922:data <=32'h00400014;14'd3923:data <=32'h003A0008;
14'd3924:data <=32'h0031FFFE;14'd3925:data <=32'h0028FFF9;14'd3926:data <=32'h001FFFF6;
14'd3927:data <=32'h0018FFF6;14'd3928:data <=32'h0010FFF7;14'd3929:data <=32'h000AFFFB;
14'd3930:data <=32'h00060000;14'd3931:data <=32'h00040007;14'd3932:data <=32'h0006000D;
14'd3933:data <=32'h000A0013;14'd3934:data <=32'h00110017;14'd3935:data <=32'h00190017;
14'd3936:data <=32'h00210013;14'd3937:data <=32'h0027000D;14'd3938:data <=32'h00290005;
14'd3939:data <=32'h0028FFFD;14'd3940:data <=32'h0025FFF6;14'd3941:data <=32'h001FFFF2;
14'd3942:data <=32'h001AFFF1;14'd3943:data <=32'h0016FFF3;14'd3944:data <=32'h0014FFF5;
14'd3945:data <=32'h0014FFF8;14'd3946:data <=32'h0016FFFB;14'd3947:data <=32'h0019FFFB;
14'd3948:data <=32'h001DFFFB;14'd3949:data <=32'h0020FFF8;14'd3950:data <=32'h0024FFF5;
14'd3951:data <=32'h0027FFF0;14'd3952:data <=32'h0029FFEB;14'd3953:data <=32'h002BFFE3;
14'd3954:data <=32'h002CFFDB;14'd3955:data <=32'h002AFFD1;14'd3956:data <=32'h0025FFC6;
14'd3957:data <=32'h001CFFBD;14'd3958:data <=32'h0011FFB7;14'd3959:data <=32'h0005FFB4;
14'd3960:data <=32'hFFF9FFB3;14'd3961:data <=32'hFFEFFFB6;14'd3962:data <=32'hFFE6FFBA;
14'd3963:data <=32'hFFE0FFBE;14'd3964:data <=32'hFFDBFFC1;14'd3965:data <=32'hFFD6FFC3;
14'd3966:data <=32'hFFCFFFC4;14'd3967:data <=32'hFFC6FFC6;14'd3968:data <=32'hFF98FFE1;
14'd3969:data <=32'hFF91FFF2;14'd3970:data <=32'hFF94FFFD;14'd3971:data <=32'hFFACFFCF;
14'd3972:data <=32'hFFA8FFC0;14'd3973:data <=32'hFF9AFFCE;14'd3974:data <=32'hFF8EFFDF;
14'd3975:data <=32'hFF86FFF3;14'd3976:data <=32'hFF820009;14'd3977:data <=32'hFF830022;
14'd3978:data <=32'hFF8A003A;14'd3979:data <=32'hFF970052;14'd3980:data <=32'hFFAB0065;
14'd3981:data <=32'hFFC40072;14'd3982:data <=32'hFFE00078;14'd3983:data <=32'hFFFB0076;
14'd3984:data <=32'h0013006C;14'd3985:data <=32'h0026005D;14'd3986:data <=32'h0032004B;
14'd3987:data <=32'h00380039;14'd3988:data <=32'h003A0028;14'd3989:data <=32'h00380018;
14'd3990:data <=32'h0033000C;14'd3991:data <=32'h002B0001;14'd3992:data <=32'h0023FFFA;
14'd3993:data <=32'h0019FFF5;14'd3994:data <=32'h000EFFF4;14'd3995:data <=32'h0004FFF6;
14'd3996:data <=32'hFFFCFFFB;14'd3997:data <=32'hFFF70003;14'd3998:data <=32'hFFF5000C;
14'd3999:data <=32'hFFF70014;14'd4000:data <=32'hFFFC0019;14'd4001:data <=32'h0001001D;
14'd4002:data <=32'h0006001F;14'd4003:data <=32'h000B001F;14'd4004:data <=32'h000F001F;
14'd4005:data <=32'h0012001F;14'd4006:data <=32'h0015001F;14'd4007:data <=32'h00190020;
14'd4008:data <=32'h001F0021;14'd4009:data <=32'h00270020;14'd4010:data <=32'h002F001C;
14'd4011:data <=32'h00360016;14'd4012:data <=32'h003C000E;14'd4013:data <=32'h003F0004;
14'd4014:data <=32'h0040FFF9;14'd4015:data <=32'h003EFFF0;14'd4016:data <=32'h003BFFE7;
14'd4017:data <=32'h0036FFDF;14'd4018:data <=32'h0030FFD9;14'd4019:data <=32'h002AFFD4;
14'd4020:data <=32'h0022FFD0;14'd4021:data <=32'h001AFFCE;14'd4022:data <=32'h0012FFCD;
14'd4023:data <=32'h000BFFD0;14'd4024:data <=32'h0005FFD4;14'd4025:data <=32'h0003FFDA;
14'd4026:data <=32'h0004FFDF;14'd4027:data <=32'h0009FFE2;14'd4028:data <=32'h000FFFE1;
14'd4029:data <=32'h0015FFDB;14'd4030:data <=32'h0019FFD1;14'd4031:data <=32'h0017FFC5;
14'd4032:data <=32'hFFE7FFAA;14'd4033:data <=32'hFFD7FFA8;14'd4034:data <=32'hFFD0FFB1;
14'd4035:data <=32'hFFF9FFBE;14'd4036:data <=32'hFFF5FFA0;14'd4037:data <=32'hFFE3FF9F;
14'd4038:data <=32'hFFCFFFA1;14'd4039:data <=32'hFFBDFFA8;14'd4040:data <=32'hFFABFFB3;
14'd4041:data <=32'hFF9BFFC3;14'd4042:data <=32'hFF8FFFD7;14'd4043:data <=32'hFF89FFEE;
14'd4044:data <=32'hFF890007;14'd4045:data <=32'hFF90001E;14'd4046:data <=32'hFF9D0032;
14'd4047:data <=32'hFFAE0040;14'd4048:data <=32'hFFC00048;14'd4049:data <=32'hFFD1004C;
14'd4050:data <=32'hFFE1004B;14'd4051:data <=32'hFFED0048;14'd4052:data <=32'hFFF80043;
14'd4053:data <=32'h0001003E;14'd4054:data <=32'h00090039;14'd4055:data <=32'h00100032;
14'd4056:data <=32'h0015002B;14'd4057:data <=32'h00180022;14'd4058:data <=32'h00190019;
14'd4059:data <=32'h00180011;14'd4060:data <=32'h0014000B;14'd4061:data <=32'h00100005;
14'd4062:data <=32'h000B0003;14'd4063:data <=32'h00060001;14'd4064:data <=32'h00010001;
14'd4065:data <=32'hFFFD0001;14'd4066:data <=32'hFFF80002;14'd4067:data <=32'hFFF20004;
14'd4068:data <=32'hFFEC0009;14'd4069:data <=32'hFFE70010;14'd4070:data <=32'hFFE4001A;
14'd4071:data <=32'hFFE50027;14'd4072:data <=32'hFFEA0033;14'd4073:data <=32'hFFF4003E;
14'd4074:data <=32'h00020047;14'd4075:data <=32'h0012004A;14'd4076:data <=32'h00230049;
14'd4077:data <=32'h00330043;14'd4078:data <=32'h00410039;14'd4079:data <=32'h004B002B;
14'd4080:data <=32'h0052001D;14'd4081:data <=32'h0055000D;14'd4082:data <=32'h0054FFFF;
14'd4083:data <=32'h0051FFF1;14'd4084:data <=32'h004BFFE4;14'd4085:data <=32'h0042FFDA;
14'd4086:data <=32'h0037FFD2;14'd4087:data <=32'h002BFFCF;14'd4088:data <=32'h001FFFD0;
14'd4089:data <=32'h0016FFD4;14'd4090:data <=32'h0011FFDB;14'd4091:data <=32'h0010FFE2;
14'd4092:data <=32'h0014FFE7;14'd4093:data <=32'h001AFFE8;14'd4094:data <=32'h0021FFE4;
14'd4095:data <=32'h0025FFDD;14'd4096:data <=32'h0029FFE0;14'd4097:data <=32'h002CFFD1;
14'd4098:data <=32'h0025FFC8;14'd4099:data <=32'h0009FFCD;14'd4100:data <=32'h000CFFB2;
14'd4101:data <=32'h0000FFB0;14'd4102:data <=32'hFFF5FFB1;14'd4103:data <=32'hFFEBFFB4;
14'd4104:data <=32'hFFE0FFB7;14'd4105:data <=32'hFFD6FFBD;14'd4106:data <=32'hFFCDFFC4;
14'd4107:data <=32'hFFC5FFCE;14'd4108:data <=32'hFFC1FFDA;14'd4109:data <=32'hFFC0FFE5;
14'd4110:data <=32'hFFC1FFF0;14'd4111:data <=32'hFFC6FFF7;14'd4112:data <=32'hFFCAFFFC;
14'd4113:data <=32'hFFCDFFFE;14'd4114:data <=32'hFFCF0000;14'd4115:data <=32'hFFCE0001;
14'd4116:data <=32'hFFCC0005;14'd4117:data <=32'hFFCB000B;14'd4118:data <=32'hFFCB0013;
14'd4119:data <=32'hFFCD001B;14'd4120:data <=32'hFFD30023;14'd4121:data <=32'hFFDB0029;
14'd4122:data <=32'hFFE3002D;14'd4123:data <=32'hFFEC002E;14'd4124:data <=32'hFFF5002D;
14'd4125:data <=32'hFFFD002B;14'd4126:data <=32'h00040026;14'd4127:data <=32'h000A0020;
14'd4128:data <=32'h000F0019;14'd4129:data <=32'h00100010;14'd4130:data <=32'h000F0006;
14'd4131:data <=32'h000AFFFD;14'd4132:data <=32'h0002FFF7;14'd4133:data <=32'hFFF6FFF3;
14'd4134:data <=32'hFFE9FFF4;14'd4135:data <=32'hFFDEFFFB;14'd4136:data <=32'hFFD50006;
14'd4137:data <=32'hFFD10014;14'd4138:data <=32'hFFD10023;14'd4139:data <=32'hFFD60032;
14'd4140:data <=32'hFFE0003D;14'd4141:data <=32'hFFEC0046;14'd4142:data <=32'hFFF9004B;
14'd4143:data <=32'h0006004D;14'd4144:data <=32'h0013004D;14'd4145:data <=32'h0020004A;
14'd4146:data <=32'h002B0045;14'd4147:data <=32'h0035003E;14'd4148:data <=32'h003F0036;
14'd4149:data <=32'h0046002C;14'd4150:data <=32'h004A0021;14'd4151:data <=32'h004C0016;
14'd4152:data <=32'h004C000C;14'd4153:data <=32'h004B0004;14'd4154:data <=32'h004AFFFD;
14'd4155:data <=32'h0049FFF8;14'd4156:data <=32'h004AFFF2;14'd4157:data <=32'h004CFFEA;
14'd4158:data <=32'h004CFFE0;14'd4159:data <=32'h004BFFD3;14'd4160:data <=32'h00160009;
14'd4161:data <=32'h00260007;14'd4162:data <=32'h0032FFFA;14'd4163:data <=32'h0032FFB8;
14'd4164:data <=32'h002CFF9B;14'd4165:data <=32'h0017FF99;14'd4166:data <=32'h0004FF9D;
14'd4167:data <=32'hFFF4FFA4;14'd4168:data <=32'hFFE7FFAE;14'd4169:data <=32'hFFDDFFB9;
14'd4170:data <=32'hFFD6FFC6;14'd4171:data <=32'hFFD2FFD3;14'd4172:data <=32'hFFD2FFE0;
14'd4173:data <=32'hFFD6FFEB;14'd4174:data <=32'hFFDDFFF4;14'd4175:data <=32'hFFE6FFF8;
14'd4176:data <=32'hFFEFFFF8;14'd4177:data <=32'hFFF7FFF3;14'd4178:data <=32'hFFFAFFEB;
14'd4179:data <=32'hFFF8FFE4;14'd4180:data <=32'hFFF2FFDD;14'd4181:data <=32'hFFE9FFDA;
14'd4182:data <=32'hFFDFFFDB;14'd4183:data <=32'hFFD6FFE0;14'd4184:data <=32'hFFCFFFE7;
14'd4185:data <=32'hFFCBFFF0;14'd4186:data <=32'hFFC9FFFA;14'd4187:data <=32'hFFCA0003;
14'd4188:data <=32'hFFCD000B;14'd4189:data <=32'hFFD10012;14'd4190:data <=32'hFFD70019;
14'd4191:data <=32'hFFDE001E;14'd4192:data <=32'hFFE70020;14'd4193:data <=32'hFFF00020;
14'd4194:data <=32'hFFF8001C;14'd4195:data <=32'hFFFD0017;14'd4196:data <=32'h0000000F;
14'd4197:data <=32'hFFFF0007;14'd4198:data <=32'hFFFB0001;14'd4199:data <=32'hFFF5FFFD;
14'd4200:data <=32'hFFEEFFFD;14'd4201:data <=32'hFFE8FFFF;14'd4202:data <=32'hFFE30003;
14'd4203:data <=32'hFFE00008;14'd4204:data <=32'hFFDF000D;14'd4205:data <=32'hFFDE0012;
14'd4206:data <=32'hFFDD0016;14'd4207:data <=32'hFFDD001A;14'd4208:data <=32'hFFDC0020;
14'd4209:data <=32'hFFDB0027;14'd4210:data <=32'hFFDC0030;14'd4211:data <=32'hFFDF0039;
14'd4212:data <=32'hFFE50043;14'd4213:data <=32'hFFED004C;14'd4214:data <=32'hFFF80054;
14'd4215:data <=32'h00050059;14'd4216:data <=32'h0013005C;14'd4217:data <=32'h0022005E;
14'd4218:data <=32'h0032005D;14'd4219:data <=32'h00440059;14'd4220:data <=32'h00570051;
14'd4221:data <=32'h00690044;14'd4222:data <=32'h00790031;14'd4223:data <=32'h00850019;
14'd4224:data <=32'h0021000A;14'd4225:data <=32'h002C000D;14'd4226:data <=32'h003E000E;
14'd4227:data <=32'h007AFFF4;14'd4228:data <=32'h007BFFC6;14'd4229:data <=32'h0068FFB3;
14'd4230:data <=32'h0053FFA5;14'd4231:data <=32'h003DFF9E;14'd4232:data <=32'h0028FF9D;
14'd4233:data <=32'h0014FF9F;14'd4234:data <=32'h0002FFA5;14'd4235:data <=32'hFFF3FFAE;
14'd4236:data <=32'hFFE8FFBB;14'd4237:data <=32'hFFE1FFC9;14'd4238:data <=32'hFFDFFFD8;
14'd4239:data <=32'hFFE2FFE4;14'd4240:data <=32'hFFE9FFEC;14'd4241:data <=32'hFFF1FFF0;
14'd4242:data <=32'hFFF8FFEF;14'd4243:data <=32'hFFFCFFEC;14'd4244:data <=32'hFFFDFFE7;
14'd4245:data <=32'hFFFBFFE3;14'd4246:data <=32'hFFF7FFE1;14'd4247:data <=32'hFFF3FFE1;
14'd4248:data <=32'hFFEFFFE2;14'd4249:data <=32'hFFECFFE5;14'd4250:data <=32'hFFEBFFE6;
14'd4251:data <=32'hFFE9FFE8;14'd4252:data <=32'hFFE8FFE9;14'd4253:data <=32'hFFE6FFEA;
14'd4254:data <=32'hFFE4FFED;14'd4255:data <=32'hFFE2FFEF;14'd4256:data <=32'hFFE1FFF3;
14'd4257:data <=32'hFFE1FFF6;14'd4258:data <=32'hFFE1FFF8;14'd4259:data <=32'hFFE1FFFB;
14'd4260:data <=32'hFFE2FFFC;14'd4261:data <=32'hFFE2FFFD;14'd4262:data <=32'hFFE1FFFF;
14'd4263:data <=32'hFFE00001;14'd4264:data <=32'hFFDF0004;14'd4265:data <=32'hFFE00009;
14'd4266:data <=32'hFFE2000D;14'd4267:data <=32'hFFE6000F;14'd4268:data <=32'hFFEB0010;
14'd4269:data <=32'hFFF0000E;14'd4270:data <=32'hFFF30009;14'd4271:data <=32'hFFF20003;
14'd4272:data <=32'hFFEDFFFD;14'd4273:data <=32'hFFE6FFFA;14'd4274:data <=32'hFFDCFFF9;
14'd4275:data <=32'hFFD2FFFE;14'd4276:data <=32'hFFC80006;14'd4277:data <=32'hFFC00011;
14'd4278:data <=32'hFFBC0020;14'd4279:data <=32'hFFBB0030;14'd4280:data <=32'hFFBE0041;
14'd4281:data <=32'hFFC60052;14'd4282:data <=32'hFFD20063;14'd4283:data <=32'hFFE30073;
14'd4284:data <=32'hFFF9007E;14'd4285:data <=32'h00130084;14'd4286:data <=32'h002F0083;
14'd4287:data <=32'h004C0079;14'd4288:data <=32'h00280049;14'd4289:data <=32'h003B004B;
14'd4290:data <=32'h0047004D;14'd4291:data <=32'h0053005B;14'd4292:data <=32'h006A0031;
14'd4293:data <=32'h006C001E;14'd4294:data <=32'h006A000D;14'd4295:data <=32'h0066FFFD;
14'd4296:data <=32'h0060FFF0;14'd4297:data <=32'h0059FFE4;14'd4298:data <=32'h0051FFD9;
14'd4299:data <=32'h0047FFD0;14'd4300:data <=32'h003CFFCA;14'd4301:data <=32'h0031FFC7;
14'd4302:data <=32'h0027FFC5;14'd4303:data <=32'h001FFFC6;14'd4304:data <=32'h0018FFC7;
14'd4305:data <=32'h0013FFC7;14'd4306:data <=32'h000DFFC7;14'd4307:data <=32'h0006FFC7;
14'd4308:data <=32'hFFFEFFC7;14'd4309:data <=32'hFFF5FFCA;14'd4310:data <=32'hFFECFFCF;
14'd4311:data <=32'hFFE6FFD8;14'd4312:data <=32'hFFE3FFE2;14'd4313:data <=32'hFFE3FFEC;
14'd4314:data <=32'hFFE7FFF5;14'd4315:data <=32'hFFEEFFFB;14'd4316:data <=32'hFFF5FFFD;
14'd4317:data <=32'hFFFCFFFD;14'd4318:data <=32'h0002FFFA;14'd4319:data <=32'h0006FFF5;
14'd4320:data <=32'h0008FFF0;14'd4321:data <=32'h0008FFEA;14'd4322:data <=32'h0006FFE4;
14'd4323:data <=32'h0003FFDF;14'd4324:data <=32'hFFFEFFDA;14'd4325:data <=32'hFFF7FFD6;
14'd4326:data <=32'hFFEEFFD5;14'd4327:data <=32'hFFE5FFD6;14'd4328:data <=32'hFFDCFFDA;
14'd4329:data <=32'hFFD5FFE2;14'd4330:data <=32'hFFD1FFEB;14'd4331:data <=32'hFFD0FFF5;
14'd4332:data <=32'hFFD4FFFD;14'd4333:data <=32'hFFD90003;14'd4334:data <=32'hFFDF0005;
14'd4335:data <=32'hFFE40003;14'd4336:data <=32'hFFE7FFFF;14'd4337:data <=32'hFFE6FFFB;
14'd4338:data <=32'hFFE3FFF7;14'd4339:data <=32'hFFDDFFF5;14'd4340:data <=32'hFFD5FFF6;
14'd4341:data <=32'hFFCDFFFA;14'd4342:data <=32'hFFC70000;14'd4343:data <=32'hFFC10008;
14'd4344:data <=32'hFFBD0012;14'd4345:data <=32'hFFBA001E;14'd4346:data <=32'hFFBA002B;
14'd4347:data <=32'hFFBD003A;14'd4348:data <=32'hFFC40049;14'd4349:data <=32'hFFCF0057;
14'd4350:data <=32'hFFE00062;14'd4351:data <=32'hFFF20068;14'd4352:data <=32'hFFD0006C;
14'd4353:data <=32'hFFE60081;14'd4354:data <=32'hFFFB0085;14'd4355:data <=32'hFFFD0058;
14'd4356:data <=32'h0012003F;14'd4357:data <=32'h0015003D;14'd4358:data <=32'h0018003C;
14'd4359:data <=32'h001B003D;14'd4360:data <=32'h0022003E;14'd4361:data <=32'h002B003D;
14'd4362:data <=32'h0035003A;14'd4363:data <=32'h003F0035;14'd4364:data <=32'h0049002C;
14'd4365:data <=32'h00500022;14'd4366:data <=32'h00560016;14'd4367:data <=32'h005A000A;
14'd4368:data <=32'h005CFFFC;14'd4369:data <=32'h005CFFEC;14'd4370:data <=32'h0058FFDB;
14'd4371:data <=32'h004FFFCB;14'd4372:data <=32'h0042FFBD;14'd4373:data <=32'h0030FFB3;
14'd4374:data <=32'h001DFFAE;14'd4375:data <=32'h0009FFB1;14'd4376:data <=32'hFFF6FFB8;
14'd4377:data <=32'hFFE9FFC5;14'd4378:data <=32'hFFE1FFD4;14'd4379:data <=32'hFFDFFFE2;
14'd4380:data <=32'hFFE1FFF0;14'd4381:data <=32'hFFE6FFFB;14'd4382:data <=32'hFFEE0002;
14'd4383:data <=32'hFFF70007;14'd4384:data <=32'h00000009;14'd4385:data <=32'h00090008;
14'd4386:data <=32'h00110005;14'd4387:data <=32'h0019FFFF;14'd4388:data <=32'h001EFFF7;
14'd4389:data <=32'h0020FFED;14'd4390:data <=32'h001FFFE3;14'd4391:data <=32'h001BFFD9;
14'd4392:data <=32'h0014FFD1;14'd4393:data <=32'h000BFFCC;14'd4394:data <=32'h0002FFCA;
14'd4395:data <=32'hFFFAFFCA;14'd4396:data <=32'hFFF3FFCC;14'd4397:data <=32'hFFEEFFCD;
14'd4398:data <=32'hFFEAFFCE;14'd4399:data <=32'hFFE5FFCF;14'd4400:data <=32'hFFDFFFCE;
14'd4401:data <=32'hFFD7FFCF;14'd4402:data <=32'hFFCEFFD1;14'd4403:data <=32'hFFC5FFD6;
14'd4404:data <=32'hFFBBFFDE;14'd4405:data <=32'hFFB5FFE9;14'd4406:data <=32'hFFB0FFF5;
14'd4407:data <=32'hFFAF0001;14'd4408:data <=32'hFFB0000E;14'd4409:data <=32'hFFB30019;
14'd4410:data <=32'hFFB80024;14'd4411:data <=32'hFFBE002D;14'd4412:data <=32'hFFC60035;
14'd4413:data <=32'hFFD0003C;14'd4414:data <=32'hFFDB0041;14'd4415:data <=32'hFFE70042;
14'd4416:data <=32'hFF970023;14'd4417:data <=32'hFF980041;14'd4418:data <=32'hFFAA0057;
14'd4419:data <=32'hFFEF003A;14'd4420:data <=32'hFFFE001E;14'd4421:data <=32'hFFF80019;
14'd4422:data <=32'hFFF0001A;14'd4423:data <=32'hFFE9001F;14'd4424:data <=32'hFFE60028;
14'd4425:data <=32'hFFE70033;14'd4426:data <=32'hFFED003D;14'd4427:data <=32'hFFF50046;
14'd4428:data <=32'h0001004D;14'd4429:data <=32'h000F0050;14'd4430:data <=32'h001D0050;
14'd4431:data <=32'h002C004E;14'd4432:data <=32'h003C0048;14'd4433:data <=32'h004A003D;
14'd4434:data <=32'h0056002E;14'd4435:data <=32'h005E001C;14'd4436:data <=32'h00610008;
14'd4437:data <=32'h005DFFF3;14'd4438:data <=32'h0054FFE1;14'd4439:data <=32'h0046FFD4;
14'd4440:data <=32'h0036FFCB;14'd4441:data <=32'h0026FFC8;14'd4442:data <=32'h0017FFCA;
14'd4443:data <=32'h000CFFCF;14'd4444:data <=32'h0003FFD5;14'd4445:data <=32'hFFFDFFDC;
14'd4446:data <=32'hFFF9FFE3;14'd4447:data <=32'hFFF6FFEA;14'd4448:data <=32'hFFF5FFF1;
14'd4449:data <=32'hFFF6FFF9;14'd4450:data <=32'hFFF80000;14'd4451:data <=32'hFFFD0006;
14'd4452:data <=32'h0004000A;14'd4453:data <=32'h000C000C;14'd4454:data <=32'h0014000C;
14'd4455:data <=32'h001C0008;14'd4456:data <=32'h00220004;14'd4457:data <=32'h0028FFFE;
14'd4458:data <=32'h002CFFF6;14'd4459:data <=32'h002FFFEE;14'd4460:data <=32'h0032FFE5;
14'd4461:data <=32'h0033FFDA;14'd4462:data <=32'h0032FFCE;14'd4463:data <=32'h002EFFBF;
14'd4464:data <=32'h0025FFB1;14'd4465:data <=32'h0018FFA4;14'd4466:data <=32'h0006FF99;
14'd4467:data <=32'hFFF1FF94;14'd4468:data <=32'hFFD9FF96;14'd4469:data <=32'hFFC3FF9D;
14'd4470:data <=32'hFFAFFFAA;14'd4471:data <=32'hFFA0FFBC;14'd4472:data <=32'hFF96FFD0;
14'd4473:data <=32'hFF91FFE5;14'd4474:data <=32'hFF91FFFA;14'd4475:data <=32'hFF95000D;
14'd4476:data <=32'hFF9D001F;14'd4477:data <=32'hFFA9002E;14'd4478:data <=32'hFFB8003A;
14'd4479:data <=32'hFFC80041;14'd4480:data <=32'hFFB8FFF6;14'd4481:data <=32'hFFAE0004;
14'd4482:data <=32'hFFAB001B;14'd4483:data <=32'hFFCE0041;14'd4484:data <=32'hFFE70027;
14'd4485:data <=32'hFFE80021;14'd4486:data <=32'hFFE6001E;14'd4487:data <=32'hFFE3001E;
14'd4488:data <=32'hFFE00021;14'd4489:data <=32'hFFDF0027;14'd4490:data <=32'hFFE1002E;
14'd4491:data <=32'hFFE50034;14'd4492:data <=32'hFFEB0038;14'd4493:data <=32'hFFF2003C;
14'd4494:data <=32'hFFF9003F;14'd4495:data <=32'h00010041;14'd4496:data <=32'h000A0041;
14'd4497:data <=32'h00140040;14'd4498:data <=32'h001E003D;14'd4499:data <=32'h00270036;
14'd4500:data <=32'h002F002D;14'd4501:data <=32'h00330024;14'd4502:data <=32'h00340019;
14'd4503:data <=32'h00320010;14'd4504:data <=32'h002E0009;14'd4505:data <=32'h002A0005;
14'd4506:data <=32'h00270002;14'd4507:data <=32'h00250001;14'd4508:data <=32'h0024FFFE;
14'd4509:data <=32'h0024FFFC;14'd4510:data <=32'h0023FFF8;14'd4511:data <=32'h0020FFF3;
14'd4512:data <=32'h001CFFEF;14'd4513:data <=32'h0016FFEC;14'd4514:data <=32'h000FFFEC;
14'd4515:data <=32'h0009FFEE;14'd4516:data <=32'h0004FFF3;14'd4517:data <=32'h0001FFF9;
14'd4518:data <=32'h0000FFFF;14'd4519:data <=32'h00010005;14'd4520:data <=32'h0004000C;
14'd4521:data <=32'h00090011;14'd4522:data <=32'h00110016;14'd4523:data <=32'h001A0019;
14'd4524:data <=32'h00260019;14'd4525:data <=32'h00330016;14'd4526:data <=32'h0040000D;
14'd4527:data <=32'h004C0000;14'd4528:data <=32'h0054FFEE;14'd4529:data <=32'h0057FFD9;
14'd4530:data <=32'h0052FFC3;14'd4531:data <=32'h0048FFAE;14'd4532:data <=32'h0037FF9C;
14'd4533:data <=32'h0022FF91;14'd4534:data <=32'h000BFF8B;14'd4535:data <=32'hFFF4FF8B;
14'd4536:data <=32'hFFDFFF90;14'd4537:data <=32'hFFCDFF99;14'd4538:data <=32'hFFBDFFA5;
14'd4539:data <=32'hFFB0FFB3;14'd4540:data <=32'hFFA6FFC3;14'd4541:data <=32'hFFA0FFD4;
14'd4542:data <=32'hFF9FFFE6;14'd4543:data <=32'hFFA1FFF6;14'd4544:data <=32'hFFB6FFF6;
14'd4545:data <=32'hFFB4FFFE;14'd4546:data <=32'hFFAE0004;14'd4547:data <=32'hFF9AFFFD;
14'd4548:data <=32'hFFACFFF2;14'd4549:data <=32'hFFAAFFFB;14'd4550:data <=32'hFFA70005;
14'd4551:data <=32'hFFA60011;14'd4552:data <=32'hFFA80020;14'd4553:data <=32'hFFAD002F;
14'd4554:data <=32'hFFB8003D;14'd4555:data <=32'hFFC50047;14'd4556:data <=32'hFFD5004D;
14'd4557:data <=32'hFFE50050;14'd4558:data <=32'hFFF3004D;14'd4559:data <=32'h00000048;
14'd4560:data <=32'h000A0042;14'd4561:data <=32'h0012003B;14'd4562:data <=32'h00180032;
14'd4563:data <=32'h001C0029;14'd4564:data <=32'h001E001F;14'd4565:data <=32'h001C0016;
14'd4566:data <=32'h0017000E;14'd4567:data <=32'h00110008;14'd4568:data <=32'h00090007;
14'd4569:data <=32'h0002000A;14'd4570:data <=32'hFFFE000F;14'd4571:data <=32'hFFFD0016;
14'd4572:data <=32'h0000001D;14'd4573:data <=32'h00060022;14'd4574:data <=32'h000E0023;
14'd4575:data <=32'h00150021;14'd4576:data <=32'h001B001D;14'd4577:data <=32'h001F0017;
14'd4578:data <=32'h00200010;14'd4579:data <=32'h001F000B;14'd4580:data <=32'h001D0007;
14'd4581:data <=32'h001A0004;14'd4582:data <=32'h00170002;14'd4583:data <=32'h00140002;
14'd4584:data <=32'h00110003;14'd4585:data <=32'h000E0006;14'd4586:data <=32'h000D000A;
14'd4587:data <=32'h000D000F;14'd4588:data <=32'h00110014;14'd4589:data <=32'h00170019;
14'd4590:data <=32'h0020001C;14'd4591:data <=32'h002B001B;14'd4592:data <=32'h00360016;
14'd4593:data <=32'h0040000D;14'd4594:data <=32'h00470000;14'd4595:data <=32'h004AFFF3;
14'd4596:data <=32'h0049FFE5;14'd4597:data <=32'h0044FFD8;14'd4598:data <=32'h003DFFCE;
14'd4599:data <=32'h0036FFC6;14'd4600:data <=32'h002EFFC0;14'd4601:data <=32'h0027FFBB;
14'd4602:data <=32'h0020FFB5;14'd4603:data <=32'h0018FFB0;14'd4604:data <=32'h000EFFAC;
14'd4605:data <=32'h0003FFA8;14'd4606:data <=32'hFFF8FFA7;14'd4607:data <=32'hFFEBFFA7;
14'd4608:data <=32'hFFBBFFBC;14'd4609:data <=32'hFFB3FFC7;14'd4610:data <=32'hFFB4FFCD;
14'd4611:data <=32'hFFD8FFA4;14'd4612:data <=32'hFFD9FF91;14'd4613:data <=32'hFFC3FF95;
14'd4614:data <=32'hFFADFF9E;14'd4615:data <=32'hFF98FFAD;14'd4616:data <=32'hFF87FFC3;
14'd4617:data <=32'hFF7DFFDD;14'd4618:data <=32'hFF7AFFFA;14'd4619:data <=32'hFF800015;
14'd4620:data <=32'hFF8C002D;14'd4621:data <=32'hFF9D0041;14'd4622:data <=32'hFFB1004E;
14'd4623:data <=32'hFFC50055;14'd4624:data <=32'hFFDA0057;14'd4625:data <=32'hFFED0055;
14'd4626:data <=32'hFFFE004F;14'd4627:data <=32'h000C0045;14'd4628:data <=32'h00180038;
14'd4629:data <=32'h001E002A;14'd4630:data <=32'h0020001B;14'd4631:data <=32'h001C000D;
14'd4632:data <=32'h00140003;14'd4633:data <=32'h000AFFFD;14'd4634:data <=32'h0000FFFC;
14'd4635:data <=32'hFFF7FFFF;14'd4636:data <=32'hFFF10005;14'd4637:data <=32'hFFEE000B;
14'd4638:data <=32'hFFEE0012;14'd4639:data <=32'hFFF00017;14'd4640:data <=32'hFFF3001A;
14'd4641:data <=32'hFFF5001C;14'd4642:data <=32'hFFF7001E;14'd4643:data <=32'hFFFA0020;
14'd4644:data <=32'hFFFC0023;14'd4645:data <=32'hFFFF0025;14'd4646:data <=32'h00030027;
14'd4647:data <=32'h00080029;14'd4648:data <=32'h000D0029;14'd4649:data <=32'h00130029;
14'd4650:data <=32'h00180028;14'd4651:data <=32'h001C0025;14'd4652:data <=32'h00200023;
14'd4653:data <=32'h00240021;14'd4654:data <=32'h0029001E;14'd4655:data <=32'h002E001A;
14'd4656:data <=32'h00330014;14'd4657:data <=32'h0036000C;14'd4658:data <=32'h00370005;
14'd4659:data <=32'h0035FFFC;14'd4660:data <=32'h0031FFF5;14'd4661:data <=32'h002BFFF2;
14'd4662:data <=32'h0025FFF1;14'd4663:data <=32'h0022FFF3;14'd4664:data <=32'h0021FFF7;
14'd4665:data <=32'h0024FFFA;14'd4666:data <=32'h002AFFFB;14'd4667:data <=32'h0031FFF8;
14'd4668:data <=32'h0039FFF2;14'd4669:data <=32'h003FFFE9;14'd4670:data <=32'h0042FFDC;
14'd4671:data <=32'h0043FFCF;14'd4672:data <=32'h0014FFAB;14'd4673:data <=32'h000BFFA6;
14'd4674:data <=32'h0006FFAB;14'd4675:data <=32'h0031FFC0;14'd4676:data <=32'h0039FF9D;
14'd4677:data <=32'h0027FF8E;14'd4678:data <=32'h0010FF83;14'd4679:data <=32'hFFF6FF7E;
14'd4680:data <=32'hFFDBFF81;14'd4681:data <=32'hFFC1FF8C;14'd4682:data <=32'hFFACFF9E;
14'd4683:data <=32'hFF9DFFB3;14'd4684:data <=32'hFF96FFCB;14'd4685:data <=32'hFF94FFE1;
14'd4686:data <=32'hFF96FFF5;14'd4687:data <=32'hFF9C0007;14'd4688:data <=32'hFFA50016;
14'd4689:data <=32'hFFB00022;14'd4690:data <=32'hFFBC002C;14'd4691:data <=32'hFFC90033;
14'd4692:data <=32'hFFD70036;14'd4693:data <=32'hFFE50036;14'd4694:data <=32'hFFF00032;
14'd4695:data <=32'hFFFA002B;14'd4696:data <=32'h00000023;14'd4697:data <=32'h0002001C;
14'd4698:data <=32'h00030016;14'd4699:data <=32'h00020012;14'd4700:data <=32'h0001000F;
14'd4701:data <=32'h0001000C;14'd4702:data <=32'h00010008;14'd4703:data <=32'h00000005;
14'd4704:data <=32'hFFFD0000;14'd4705:data <=32'hFFF8FFFC;14'd4706:data <=32'hFFF1FFFA;
14'd4707:data <=32'hFFE9FFFB;14'd4708:data <=32'hFFE0FFFF;14'd4709:data <=32'hFFD90006;
14'd4710:data <=32'hFFD50010;14'd4711:data <=32'hFFD4001C;14'd4712:data <=32'hFFD60028;
14'd4713:data <=32'hFFDB0033;14'd4714:data <=32'hFFE4003C;14'd4715:data <=32'hFFEE0044;
14'd4716:data <=32'hFFFA0049;14'd4717:data <=32'h0007004B;14'd4718:data <=32'h0015004B;
14'd4719:data <=32'h00220047;14'd4720:data <=32'h002F003F;14'd4721:data <=32'h003A0035;
14'd4722:data <=32'h00400027;14'd4723:data <=32'h00430019;14'd4724:data <=32'h0040000B;
14'd4725:data <=32'h003A0001;14'd4726:data <=32'h0031FFFA;14'd4727:data <=32'h0028FFF8;
14'd4728:data <=32'h0020FFFB;14'd4729:data <=32'h001C0000;14'd4730:data <=32'h001D0006;
14'd4731:data <=32'h0021000B;14'd4732:data <=32'h0028000D;14'd4733:data <=32'h0030000C;
14'd4734:data <=32'h00390008;14'd4735:data <=32'h00410002;14'd4736:data <=32'h003CFFFE;
14'd4737:data <=32'h0047FFF6;14'd4738:data <=32'h0048FFED;14'd4739:data <=32'h0034FFEE;
14'd4740:data <=32'h0047FFD1;14'd4741:data <=32'h0041FFC4;14'd4742:data <=32'h0037FFB8;
14'd4743:data <=32'h002AFFAD;14'd4744:data <=32'h001BFFA8;14'd4745:data <=32'h000BFFA7;
14'd4746:data <=32'hFFFCFFAB;14'd4747:data <=32'hFFF0FFB1;14'd4748:data <=32'hFFE7FFB9;
14'd4749:data <=32'hFFE2FFC0;14'd4750:data <=32'hFFDEFFC7;14'd4751:data <=32'hFFDBFFCB;
14'd4752:data <=32'hFFD8FFD0;14'd4753:data <=32'hFFD3FFD4;14'd4754:data <=32'hFFCEFFDA;
14'd4755:data <=32'hFFCAFFE0;14'd4756:data <=32'hFFC7FFE8;14'd4757:data <=32'hFFC7FFF0;
14'd4758:data <=32'hFFC7FFF8;14'd4759:data <=32'hFFC8FFFF;14'd4760:data <=32'hFFCA0006;
14'd4761:data <=32'hFFCD000D;14'd4762:data <=32'hFFD10013;14'd4763:data <=32'hFFD6001A;
14'd4764:data <=32'hFFDE0020;14'd4765:data <=32'hFFE80023;14'd4766:data <=32'hFFF30023;
14'd4767:data <=32'hFFFE001F;14'd4768:data <=32'h00070017;14'd4769:data <=32'h000C000C;
14'd4770:data <=32'h000C0000;14'd4771:data <=32'h0007FFF5;14'd4772:data <=32'hFFFFFFEC;
14'd4773:data <=32'hFFF3FFE7;14'd4774:data <=32'hFFE7FFE7;14'd4775:data <=32'hFFDBFFEB;
14'd4776:data <=32'hFFD0FFF2;14'd4777:data <=32'hFFC9FFFC;14'd4778:data <=32'hFFC40008;
14'd4779:data <=32'hFFC20015;14'd4780:data <=32'hFFC30021;14'd4781:data <=32'hFFC7002F;
14'd4782:data <=32'hFFCE003B;14'd4783:data <=32'hFFD80045;14'd4784:data <=32'hFFE5004E;
14'd4785:data <=32'hFFF40051;14'd4786:data <=32'h00020051;14'd4787:data <=32'h000F004E;
14'd4788:data <=32'h00190047;14'd4789:data <=32'h0020003F;14'd4790:data <=32'h00240039;
14'd4791:data <=32'h00260033;14'd4792:data <=32'h00290030;14'd4793:data <=32'h002C002F;
14'd4794:data <=32'h0031002E;14'd4795:data <=32'h0037002B;14'd4796:data <=32'h003F0026;
14'd4797:data <=32'h0046001F;14'd4798:data <=32'h004C0015;14'd4799:data <=32'h0050000B;
14'd4800:data <=32'h000B0026;14'd4801:data <=32'h001C0030;14'd4802:data <=32'h0030002C;
14'd4803:data <=32'h0047FFF2;14'd4804:data <=32'h0054FFD6;14'd4805:data <=32'h004AFFCA;
14'd4806:data <=32'h003CFFC1;14'd4807:data <=32'h002EFFBC;14'd4808:data <=32'h001EFFBB;
14'd4809:data <=32'h000FFFBE;14'd4810:data <=32'h0004FFC6;14'd4811:data <=32'hFFFDFFD0;
14'd4812:data <=32'hFFFBFFDB;14'd4813:data <=32'hFFFDFFE3;14'd4814:data <=32'h0003FFE8;
14'd4815:data <=32'h0009FFE8;14'd4816:data <=32'h000EFFE4;14'd4817:data <=32'h0010FFDE;
14'd4818:data <=32'h000FFFD7;14'd4819:data <=32'h000AFFD1;14'd4820:data <=32'h0004FFCC;
14'd4821:data <=32'hFFFCFFC9;14'd4822:data <=32'hFFF4FFC8;14'd4823:data <=32'hFFEBFFC8;
14'd4824:data <=32'hFFE1FFCB;14'd4825:data <=32'hFFD7FFD0;14'd4826:data <=32'hFFCFFFD8;
14'd4827:data <=32'hFFC9FFE3;14'd4828:data <=32'hFFC5FFF0;14'd4829:data <=32'hFFC7FFFD;
14'd4830:data <=32'hFFCD0009;14'd4831:data <=32'hFFD70011;14'd4832:data <=32'hFFE20016;
14'd4833:data <=32'hFFED0016;14'd4834:data <=32'hFFF60012;14'd4835:data <=32'hFFFD000B;
14'd4836:data <=32'h00000003;14'd4837:data <=32'hFFFFFFFC;14'd4838:data <=32'hFFFDFFF5;
14'd4839:data <=32'hFFF8FFF1;14'd4840:data <=32'hFFF3FFEE;14'd4841:data <=32'hFFEEFFEC;
14'd4842:data <=32'hFFE8FFEB;14'd4843:data <=32'hFFE1FFEB;14'd4844:data <=32'hFFDBFFED;
14'd4845:data <=32'hFFD4FFF0;14'd4846:data <=32'hFFCDFFF5;14'd4847:data <=32'hFFC7FFFD;
14'd4848:data <=32'hFFC20005;14'd4849:data <=32'hFFC0000F;14'd4850:data <=32'hFFC00019;
14'd4851:data <=32'hFFC10023;14'd4852:data <=32'hFFC3002D;14'd4853:data <=32'hFFC60036;
14'd4854:data <=32'hFFC90041;14'd4855:data <=32'hFFCF004C;14'd4856:data <=32'hFFD70059;
14'd4857:data <=32'hFFE40065;14'd4858:data <=32'hFFF40070;14'd4859:data <=32'h000A0076;
14'd4860:data <=32'h00210076;14'd4861:data <=32'h00390071;14'd4862:data <=32'h004E0064;
14'd4863:data <=32'h00600053;14'd4864:data <=32'h0004001E;14'd4865:data <=32'h0009002B;
14'd4866:data <=32'h001A003B;14'd4867:data <=32'h00620038;14'd4868:data <=32'h007B0012;
14'd4869:data <=32'h0077FFFA;14'd4870:data <=32'h006DFFE5;14'd4871:data <=32'h005FFFD4;
14'd4872:data <=32'h004DFFC7;14'd4873:data <=32'h0039FFC1;14'd4874:data <=32'h0026FFC1;
14'd4875:data <=32'h0016FFC6;14'd4876:data <=32'h000BFFD0;14'd4877:data <=32'h0005FFDB;
14'd4878:data <=32'h0005FFE5;14'd4879:data <=32'h0008FFEC;14'd4880:data <=32'h000DFFEF;
14'd4881:data <=32'h0011FFEF;14'd4882:data <=32'h0015FFED;14'd4883:data <=32'h0016FFE9;
14'd4884:data <=32'h0016FFE5;14'd4885:data <=32'h0015FFE2;14'd4886:data <=32'h0013FFDE;
14'd4887:data <=32'h0011FFDA;14'd4888:data <=32'h000DFFD6;14'd4889:data <=32'h0007FFD3;
14'd4890:data <=32'h0001FFD1;14'd4891:data <=32'hFFF9FFD1;14'd4892:data <=32'hFFF1FFD4;
14'd4893:data <=32'hFFECFFD9;14'd4894:data <=32'hFFE8FFDF;14'd4895:data <=32'hFFE7FFE5;
14'd4896:data <=32'hFFE8FFEA;14'd4897:data <=32'hFFEAFFED;14'd4898:data <=32'hFFECFFEF;
14'd4899:data <=32'hFFEDFFEE;14'd4900:data <=32'hFFECFFEE;14'd4901:data <=32'hFFEBFFEF;
14'd4902:data <=32'hFFE9FFF1;14'd4903:data <=32'hFFE8FFF4;14'd4904:data <=32'hFFE9FFF8;
14'd4905:data <=32'hFFEBFFFA;14'd4906:data <=32'hFFEFFFFC;14'd4907:data <=32'hFFF3FFFB;
14'd4908:data <=32'hFFF6FFF7;14'd4909:data <=32'hFFF8FFF2;14'd4910:data <=32'hFFF7FFEC;
14'd4911:data <=32'hFFF3FFE6;14'd4912:data <=32'hFFEDFFE1;14'd4913:data <=32'hFFE5FFDE;
14'd4914:data <=32'hFFDCFFDB;14'd4915:data <=32'hFFD1FFDB;14'd4916:data <=32'hFFC4FFDE;
14'd4917:data <=32'hFFB7FFE4;14'd4918:data <=32'hFFA9FFEE;14'd4919:data <=32'hFF9DFFFE;
14'd4920:data <=32'hFF940012;14'd4921:data <=32'hFF91002B;14'd4922:data <=32'hFF950046;
14'd4923:data <=32'hFFA1005F;14'd4924:data <=32'hFFB40075;14'd4925:data <=32'hFFCD0085;
14'd4926:data <=32'hFFEA008D;14'd4927:data <=32'h0007008E;14'd4928:data <=32'hFFF70047;
14'd4929:data <=32'h00000053;14'd4930:data <=32'h00050061;14'd4931:data <=32'h0012007F;
14'd4932:data <=32'h003B0066;14'd4933:data <=32'h00480057;14'd4934:data <=32'h00520047;
14'd4935:data <=32'h00580035;14'd4936:data <=32'h00590023;14'd4937:data <=32'h00570014;
14'd4938:data <=32'h00510007;14'd4939:data <=32'h0049FFFE;14'd4940:data <=32'h0042FFF8;
14'd4941:data <=32'h003DFFF5;14'd4942:data <=32'h003AFFF2;14'd4943:data <=32'h0038FFEE;
14'd4944:data <=32'h0035FFE8;14'd4945:data <=32'h0032FFE2;14'd4946:data <=32'h002CFFDC;
14'd4947:data <=32'h0025FFD8;14'd4948:data <=32'h001CFFD5;14'd4949:data <=32'h0013FFD6;
14'd4950:data <=32'h000CFFD9;14'd4951:data <=32'h0007FFDD;14'd4952:data <=32'h0003FFE1;
14'd4953:data <=32'h0002FFE6;14'd4954:data <=32'h0001FFEA;14'd4955:data <=32'h0001FFED;
14'd4956:data <=32'h0001FFF1;14'd4957:data <=32'h0003FFF3;14'd4958:data <=32'h0007FFF5;
14'd4959:data <=32'h000BFFF5;14'd4960:data <=32'h0010FFF4;14'd4961:data <=32'h0014FFEF;
14'd4962:data <=32'h0016FFE9;14'd4963:data <=32'h0015FFE1;14'd4964:data <=32'h0011FFD9;
14'd4965:data <=32'h000AFFD4;14'd4966:data <=32'h0001FFD1;14'd4967:data <=32'hFFF7FFD2;
14'd4968:data <=32'hFFEFFFD6;14'd4969:data <=32'hFFEAFFDD;14'd4970:data <=32'hFFE8FFE3;
14'd4971:data <=32'hFFE9FFEA;14'd4972:data <=32'hFFECFFEE;14'd4973:data <=32'hFFF0FFF0;
14'd4974:data <=32'hFFF3FFEF;14'd4975:data <=32'hFFF6FFED;14'd4976:data <=32'hFFF7FFE9;
14'd4977:data <=32'hFFF7FFE4;14'd4978:data <=32'hFFF5FFDF;14'd4979:data <=32'hFFF1FFD8;
14'd4980:data <=32'hFFEAFFD3;14'd4981:data <=32'hFFE0FFCF;14'd4982:data <=32'hFFD3FFCC;
14'd4983:data <=32'hFFC4FFCE;14'd4984:data <=32'hFFB5FFD5;14'd4985:data <=32'hFFA6FFE2;
14'd4986:data <=32'hFF9BFFF3;14'd4987:data <=32'hFF960008;14'd4988:data <=32'hFF97001E;
14'd4989:data <=32'hFF9D0032;14'd4990:data <=32'hFFA80043;14'd4991:data <=32'hFFB60050;
14'd4992:data <=32'hFFA20043;14'd4993:data <=32'hFFA8005C;14'd4994:data <=32'hFFB20069;
14'd4995:data <=32'hFFBB004B;14'd4996:data <=32'hFFDA0044;14'd4997:data <=32'hFFE10048;
14'd4998:data <=32'hFFE9004C;14'd4999:data <=32'hFFF20050;14'd5000:data <=32'hFFFB0051;
14'd5001:data <=32'h00040052;14'd5002:data <=32'h000D0052;14'd5003:data <=32'h00170052;
14'd5004:data <=32'h00220052;14'd5005:data <=32'h002F004F;14'd5006:data <=32'h003D004A;
14'd5007:data <=32'h004B0040;14'd5008:data <=32'h00570031;14'd5009:data <=32'h005F001F;
14'd5010:data <=32'h0061000B;14'd5011:data <=32'h005EFFF6;14'd5012:data <=32'h0055FFE4;
14'd5013:data <=32'h0047FFD7;14'd5014:data <=32'h0037FFCE;14'd5015:data <=32'h0028FFCA;
14'd5016:data <=32'h0019FFCB;14'd5017:data <=32'h000CFFCF;14'd5018:data <=32'h0001FFD5;
14'd5019:data <=32'hFFF8FFDE;14'd5020:data <=32'hFFF3FFE8;14'd5021:data <=32'hFFF1FFF3;
14'd5022:data <=32'hFFF3FFFE;14'd5023:data <=32'hFFF80008;14'd5024:data <=32'h0001000F;
14'd5025:data <=32'h000C0012;14'd5026:data <=32'h00170011;14'd5027:data <=32'h0021000B;
14'd5028:data <=32'h00280003;14'd5029:data <=32'h002BFFF9;14'd5030:data <=32'h002BFFEF;
14'd5031:data <=32'h0028FFE6;14'd5032:data <=32'h0023FFE0;14'd5033:data <=32'h001EFFDC;
14'd5034:data <=32'h001AFFD9;14'd5035:data <=32'h0016FFD7;14'd5036:data <=32'h0014FFD5;
14'd5037:data <=32'h0011FFD1;14'd5038:data <=32'h000DFFCE;14'd5039:data <=32'h0008FFCA;
14'd5040:data <=32'h0002FFC8;14'd5041:data <=32'hFFFBFFC5;14'd5042:data <=32'hFFF4FFC5;
14'd5043:data <=32'hFFEDFFC5;14'd5044:data <=32'hFFE6FFC6;14'd5045:data <=32'hFFDEFFC7;
14'd5046:data <=32'hFFD7FFC9;14'd5047:data <=32'hFFCEFFCC;14'd5048:data <=32'hFFC5FFD2;
14'd5049:data <=32'hFFBCFFDC;14'd5050:data <=32'hFFB7FFE6;14'd5051:data <=32'hFFB3FFF3;
14'd5052:data <=32'hFFB50000;14'd5053:data <=32'hFFB9000B;14'd5054:data <=32'hFFC00013;
14'd5055:data <=32'hFFC70018;14'd5056:data <=32'hFF8FFFE4;14'd5057:data <=32'hFF80FFFD;
14'd5058:data <=32'hFF820015;14'd5059:data <=32'hFFC50011;14'd5060:data <=32'hFFD90004;
14'd5061:data <=32'hFFD30004;14'd5062:data <=32'hFFCD0007;14'd5063:data <=32'hFFC7000E;
14'd5064:data <=32'hFFC30017;14'd5065:data <=32'hFFC00021;14'd5066:data <=32'hFFC0002E;
14'd5067:data <=32'hFFC2003C;14'd5068:data <=32'hFFC9004B;14'd5069:data <=32'hFFD5005A;
14'd5070:data <=32'hFFE60065;14'd5071:data <=32'hFFFB006C;14'd5072:data <=32'h0012006D;
14'd5073:data <=32'h00290066;14'd5074:data <=32'h003D0059;14'd5075:data <=32'h004B0048;
14'd5076:data <=32'h00530033;14'd5077:data <=32'h0056001F;14'd5078:data <=32'h0053000D;
14'd5079:data <=32'h004DFFFE;14'd5080:data <=32'h0044FFF1;14'd5081:data <=32'h003AFFE8;
14'd5082:data <=32'h002FFFE1;14'd5083:data <=32'h0022FFDD;14'd5084:data <=32'h0016FFDD;
14'd5085:data <=32'h000BFFDF;14'd5086:data <=32'h0001FFE5;14'd5087:data <=32'hFFFAFFEE;
14'd5088:data <=32'hFFF6FFF8;14'd5089:data <=32'hFFF70001;14'd5090:data <=32'hFFFA000A;
14'd5091:data <=32'h00000010;14'd5092:data <=32'h00060013;14'd5093:data <=32'h000C0016;
14'd5094:data <=32'h00120016;14'd5095:data <=32'h00180016;14'd5096:data <=32'h001E0016;
14'd5097:data <=32'h00250015;14'd5098:data <=32'h002D0013;14'd5099:data <=32'h0036000F;
14'd5100:data <=32'h003F0006;14'd5101:data <=32'h0047FFFB;14'd5102:data <=32'h004CFFEC;
14'd5103:data <=32'h004DFFDC;14'd5104:data <=32'h0049FFCB;14'd5105:data <=32'h0041FFBA;
14'd5106:data <=32'h0034FFAD;14'd5107:data <=32'h0025FFA2;14'd5108:data <=32'h0014FF9C;
14'd5109:data <=32'h0002FF99;14'd5110:data <=32'hFFF0FF99;14'd5111:data <=32'hFFDDFF9D;
14'd5112:data <=32'hFFCCFFA6;14'd5113:data <=32'hFFBDFFB2;14'd5114:data <=32'hFFB1FFC3;
14'd5115:data <=32'hFFABFFD5;14'd5116:data <=32'hFFAAFFE9;14'd5117:data <=32'hFFB0FFFA;
14'd5118:data <=32'hFFBA0008;14'd5119:data <=32'hFFC6000F;14'd5120:data <=32'hFFCFFFC4;
14'd5121:data <=32'hFFBEFFC7;14'd5122:data <=32'hFFAEFFD6;14'd5123:data <=32'hFFC10008;
14'd5124:data <=32'hFFDBFFFB;14'd5125:data <=32'hFFDAFFF8;14'd5126:data <=32'hFFD6FFF8;
14'd5127:data <=32'hFFD1FFF9;14'd5128:data <=32'hFFCCFFFC;14'd5129:data <=32'hFFC8FFFF;
14'd5130:data <=32'hFFC30005;14'd5131:data <=32'hFFBF000D;14'd5132:data <=32'hFFBD0018;
14'd5133:data <=32'hFFBD0025;14'd5134:data <=32'hFFC20033;14'd5135:data <=32'hFFCB003F;
14'd5136:data <=32'hFFD80049;14'd5137:data <=32'hFFE7004D;14'd5138:data <=32'hFFF6004E;
14'd5139:data <=32'h0003004A;14'd5140:data <=32'h000E0044;14'd5141:data <=32'h0016003C;
14'd5142:data <=32'h001B0035;14'd5143:data <=32'h001E002E;14'd5144:data <=32'h00210028;
14'd5145:data <=32'h00230023;14'd5146:data <=32'h0026001D;14'd5147:data <=32'h00270016;
14'd5148:data <=32'h0027000F;14'd5149:data <=32'h00250008;14'd5150:data <=32'h00210002;
14'd5151:data <=32'h001CFFFE;14'd5152:data <=32'h0018FFFB;14'd5153:data <=32'h0013FFFA;
14'd5154:data <=32'h000EFFFA;14'd5155:data <=32'h0009FFFB;14'd5156:data <=32'h0005FFFC;
14'd5157:data <=32'h0000FFFF;14'd5158:data <=32'hFFFC0004;14'd5159:data <=32'hFFF8000A;
14'd5160:data <=32'hFFF70013;14'd5161:data <=32'hFFF8001E;14'd5162:data <=32'hFFFF0029;
14'd5163:data <=32'h000A0033;14'd5164:data <=32'h00190039;14'd5165:data <=32'h002B003A;
14'd5166:data <=32'h003D0035;14'd5167:data <=32'h004E002A;14'd5168:data <=32'h005C001A;
14'd5169:data <=32'h00650007;14'd5170:data <=32'h0068FFF2;14'd5171:data <=32'h0067FFDD;
14'd5172:data <=32'h0061FFC9;14'd5173:data <=32'h0056FFB7;14'd5174:data <=32'h0049FFA7;
14'd5175:data <=32'h0037FF9A;14'd5176:data <=32'h0023FF92;14'd5177:data <=32'h000DFF8E;
14'd5178:data <=32'hFFF7FF91;14'd5179:data <=32'hFFE4FF99;14'd5180:data <=32'hFFD4FFA6;
14'd5181:data <=32'hFFCAFFB5;14'd5182:data <=32'hFFC5FFC4;14'd5183:data <=32'hFFC5FFD1;
14'd5184:data <=32'hFFDEFFD6;14'd5185:data <=32'hFFDAFFD5;14'd5186:data <=32'hFFD1FFD1;
14'd5187:data <=32'hFFB9FFC6;14'd5188:data <=32'hFFC9FFC2;14'd5189:data <=32'hFFC0FFC9;
14'd5190:data <=32'hFFB9FFD2;14'd5191:data <=32'hFFB2FFDD;14'd5192:data <=32'hFFAFFFE9;
14'd5193:data <=32'hFFAEFFF6;14'd5194:data <=32'hFFB00001;14'd5195:data <=32'hFFB3000C;
14'd5196:data <=32'hFFB70017;14'd5197:data <=32'hFFBD0020;14'd5198:data <=32'hFFC50029;
14'd5199:data <=32'hFFCF0030;14'd5200:data <=32'hFFDB0034;14'd5201:data <=32'hFFE70034;
14'd5202:data <=32'hFFF30031;14'd5203:data <=32'hFFFB002A;14'd5204:data <=32'hFFFF0021;
14'd5205:data <=32'hFFFF0019;14'd5206:data <=32'hFFFC0014;14'd5207:data <=32'hFFF70012;
14'd5208:data <=32'hFFF30013;14'd5209:data <=32'hFFF00016;14'd5210:data <=32'hFFF0001B;
14'd5211:data <=32'hFFF20020;14'd5212:data <=32'hFFF60023;14'd5213:data <=32'hFFFB0025;
14'd5214:data <=32'h00000026;14'd5215:data <=32'h00050025;14'd5216:data <=32'h000A0023;
14'd5217:data <=32'h000E0021;14'd5218:data <=32'h0012001C;14'd5219:data <=32'h00150017;
14'd5220:data <=32'h00150011;14'd5221:data <=32'h0014000B;14'd5222:data <=32'h000F0006;
14'd5223:data <=32'h00080004;14'd5224:data <=32'h00010004;14'd5225:data <=32'hFFF90009;
14'd5226:data <=32'hFFF50011;14'd5227:data <=32'hFFF3001C;14'd5228:data <=32'hFFF70027;
14'd5229:data <=32'hFFFF0031;14'd5230:data <=32'h000A0037;14'd5231:data <=32'h0017003A;
14'd5232:data <=32'h00250039;14'd5233:data <=32'h00310034;14'd5234:data <=32'h003C002D;
14'd5235:data <=32'h00450025;14'd5236:data <=32'h004C001A;14'd5237:data <=32'h0052000F;
14'd5238:data <=32'h00560003;14'd5239:data <=32'h0058FFF5;14'd5240:data <=32'h0056FFE7;
14'd5241:data <=32'h0053FFDA;14'd5242:data <=32'h004CFFCE;14'd5243:data <=32'h0044FFC5;
14'd5244:data <=32'h003AFFBD;14'd5245:data <=32'h0032FFB8;14'd5246:data <=32'h002AFFB4;
14'd5247:data <=32'h0023FFAF;14'd5248:data <=32'hFFEEFFB7;14'd5249:data <=32'hFFE9FFBB;
14'd5250:data <=32'hFFECFFBA;14'd5251:data <=32'h0015FF97;14'd5252:data <=32'h001AFF84;
14'd5253:data <=32'h0001FF7E;14'd5254:data <=32'hFFE8FF7F;14'd5255:data <=32'hFFCEFF87;
14'd5256:data <=32'hFFB9FF94;14'd5257:data <=32'hFFA8FFA6;14'd5258:data <=32'hFF9BFFBB;
14'd5259:data <=32'hFF94FFD1;14'd5260:data <=32'hFF92FFE7;14'd5261:data <=32'hFF95FFFD;
14'd5262:data <=32'hFF9C0011;14'd5263:data <=32'hFFA80023;14'd5264:data <=32'hFFB80030;
14'd5265:data <=32'hFFCB0038;14'd5266:data <=32'hFFDE003A;14'd5267:data <=32'hFFF00035;
14'd5268:data <=32'hFFFD002B;14'd5269:data <=32'h0005001F;14'd5270:data <=32'h00070013;
14'd5271:data <=32'h00040008;14'd5272:data <=32'hFFFF0001;14'd5273:data <=32'hFFF8FFFE;
14'd5274:data <=32'hFFF2FFFD;14'd5275:data <=32'hFFECFFFF;14'd5276:data <=32'hFFE90002;
14'd5277:data <=32'hFFE60005;14'd5278:data <=32'hFFE40009;14'd5279:data <=32'hFFE3000D;
14'd5280:data <=32'hFFE30012;14'd5281:data <=32'hFFE40017;14'd5282:data <=32'hFFE7001B;
14'd5283:data <=32'hFFEA001F;14'd5284:data <=32'hFFEF0021;14'd5285:data <=32'hFFF30022;
14'd5286:data <=32'hFFF70021;14'd5287:data <=32'hFFF90020;14'd5288:data <=32'hFFF9001F;
14'd5289:data <=32'hFFF90020;14'd5290:data <=32'hFFF90022;14'd5291:data <=32'hFFFA0025;
14'd5292:data <=32'hFFFD0029;14'd5293:data <=32'h0002002D;14'd5294:data <=32'h0009002E;
14'd5295:data <=32'h0010002D;14'd5296:data <=32'h0016002A;14'd5297:data <=32'h001A0025;
14'd5298:data <=32'h001C0021;14'd5299:data <=32'h001C001E;14'd5300:data <=32'h001C001D;
14'd5301:data <=32'h001C001D;14'd5302:data <=32'h001D001E;14'd5303:data <=32'h00200020;
14'd5304:data <=32'h00250021;14'd5305:data <=32'h002B0022;14'd5306:data <=32'h00320021;
14'd5307:data <=32'h003A001F;14'd5308:data <=32'h0043001C;14'd5309:data <=32'h004C0016;
14'd5310:data <=32'h0057000E;14'd5311:data <=32'h00610001;14'd5312:data <=32'h0039FFCC;
14'd5313:data <=32'h0038FFC5;14'd5314:data <=32'h0038FFC6;14'd5315:data <=32'h0060FFE1;
14'd5316:data <=32'h0075FFBF;14'd5317:data <=32'h0067FFA7;14'd5318:data <=32'h0053FF93;
14'd5319:data <=32'h003AFF85;14'd5320:data <=32'h0020FF7E;14'd5321:data <=32'h0007FF7D;
14'd5322:data <=32'hFFEFFF82;14'd5323:data <=32'hFFD9FF8B;14'd5324:data <=32'hFFC6FF99;
14'd5325:data <=32'hFFB8FFA9;14'd5326:data <=32'hFFACFFBC;14'd5327:data <=32'hFFA7FFD1;
14'd5328:data <=32'hFFA7FFE6;14'd5329:data <=32'hFFACFFF8;14'd5330:data <=32'hFFB60007;
14'd5331:data <=32'hFFC20011;14'd5332:data <=32'hFFCF0017;14'd5333:data <=32'hFFDA0018;
14'd5334:data <=32'hFFE30016;14'd5335:data <=32'hFFE90013;14'd5336:data <=32'hFFED0010;
14'd5337:data <=32'hFFF0000E;14'd5338:data <=32'hFFF3000D;14'd5339:data <=32'hFFF6000B;
14'd5340:data <=32'hFFF80008;14'd5341:data <=32'hFFFB0004;14'd5342:data <=32'hFFFBFFFF;
14'd5343:data <=32'hFFFAFFFA;14'd5344:data <=32'hFFF6FFF5;14'd5345:data <=32'hFFF1FFF2;
14'd5346:data <=32'hFFEBFFF1;14'd5347:data <=32'hFFE4FFF2;14'd5348:data <=32'hFFDEFFF5;
14'd5349:data <=32'hFFD8FFF9;14'd5350:data <=32'hFFD4FFFF;14'd5351:data <=32'hFFD00005;
14'd5352:data <=32'hFFCD000C;14'd5353:data <=32'hFFCB0016;14'd5354:data <=32'hFFCB0021;
14'd5355:data <=32'hFFCE002C;14'd5356:data <=32'hFFD60037;14'd5357:data <=32'hFFE00040;
14'd5358:data <=32'hFFEE0045;14'd5359:data <=32'hFFFC0047;14'd5360:data <=32'h00090043;
14'd5361:data <=32'h0014003B;14'd5362:data <=32'h001A0031;14'd5363:data <=32'h001C0027;
14'd5364:data <=32'h001B001F;14'd5365:data <=32'h0017001A;14'd5366:data <=32'h00120017;
14'd5367:data <=32'h000E0018;14'd5368:data <=32'h000B001B;14'd5369:data <=32'h000A001F;
14'd5370:data <=32'h000A0025;14'd5371:data <=32'h000E002B;14'd5372:data <=32'h00130032;
14'd5373:data <=32'h001C0038;14'd5374:data <=32'h0029003C;14'd5375:data <=32'h0039003D;
14'd5376:data <=32'h0036002B;14'd5377:data <=32'h0048002A;14'd5378:data <=32'h00510024;
14'd5379:data <=32'h00440022;14'd5380:data <=32'h0064000A;14'd5381:data <=32'h0065FFF7;
14'd5382:data <=32'h0061FFE5;14'd5383:data <=32'h0058FFD5;14'd5384:data <=32'h004EFFCA;
14'd5385:data <=32'h0042FFC1;14'd5386:data <=32'h0037FFBB;14'd5387:data <=32'h002CFFB7;
14'd5388:data <=32'h0022FFB3;14'd5389:data <=32'h0016FFB2;14'd5390:data <=32'h000BFFB2;
14'd5391:data <=32'hFFFFFFB4;14'd5392:data <=32'hFFF6FFB8;14'd5393:data <=32'hFFEEFFBE;
14'd5394:data <=32'hFFE8FFC4;14'd5395:data <=32'hFFE3FFCA;14'd5396:data <=32'hFFE0FFCF;
14'd5397:data <=32'hFFDCFFD3;14'd5398:data <=32'hFFD8FFD7;14'd5399:data <=32'hFFD2FFDD;
14'd5400:data <=32'hFFCEFFE5;14'd5401:data <=32'hFFCBFFEF;14'd5402:data <=32'hFFCCFFFB;
14'd5403:data <=32'hFFD00005;14'd5404:data <=32'hFFD8000E;14'd5405:data <=32'hFFE30014;
14'd5406:data <=32'hFFEE0015;14'd5407:data <=32'hFFF90012;14'd5408:data <=32'h0001000C;
14'd5409:data <=32'h00070004;14'd5410:data <=32'h0009FFFA;14'd5411:data <=32'h0008FFF1;
14'd5412:data <=32'h0004FFE8;14'd5413:data <=32'hFFFDFFE1;14'd5414:data <=32'hFFF4FFDB;
14'd5415:data <=32'hFFEAFFD8;14'd5416:data <=32'hFFDEFFD8;14'd5417:data <=32'hFFD1FFDC;
14'd5418:data <=32'hFFC4FFE3;14'd5419:data <=32'hFFBBFFEF;14'd5420:data <=32'hFFB5FFFD;
14'd5421:data <=32'hFFB3000D;14'd5422:data <=32'hFFB7001D;14'd5423:data <=32'hFFBE002A;
14'd5424:data <=32'hFFC90034;14'd5425:data <=32'hFFD40039;14'd5426:data <=32'hFFDF003B;
14'd5427:data <=32'hFFE7003A;14'd5428:data <=32'hFFED003A;14'd5429:data <=32'hFFF20038;
14'd5430:data <=32'hFFF50038;14'd5431:data <=32'hFFF90039;14'd5432:data <=32'hFFFD003A;
14'd5433:data <=32'h0002003C;14'd5434:data <=32'h0007003D;14'd5435:data <=32'h000C003D;
14'd5436:data <=32'h0012003E;14'd5437:data <=32'h0018003F;14'd5438:data <=32'h001F003F;
14'd5439:data <=32'h0028003F;14'd5440:data <=32'hFFE9003C;14'd5441:data <=32'hFFF80050;
14'd5442:data <=32'h000F0057;14'd5443:data <=32'h00380029;14'd5444:data <=32'h00550014;
14'd5445:data <=32'h00520005;14'd5446:data <=32'h004AFFF7;14'd5447:data <=32'h0040FFEE;
14'd5448:data <=32'h0036FFE9;14'd5449:data <=32'h002CFFE9;14'd5450:data <=32'h0026FFEC;
14'd5451:data <=32'h0023FFEF;14'd5452:data <=32'h0022FFF1;14'd5453:data <=32'h0024FFF2;
14'd5454:data <=32'h0026FFF1;14'd5455:data <=32'h0028FFEF;14'd5456:data <=32'h002AFFEB;
14'd5457:data <=32'h002BFFE7;14'd5458:data <=32'h002CFFE1;14'd5459:data <=32'h002BFFD9;
14'd5460:data <=32'h0029FFD0;14'd5461:data <=32'h0023FFC7;14'd5462:data <=32'h001AFFBE;
14'd5463:data <=32'h000DFFB8;14'd5464:data <=32'hFFFEFFB6;14'd5465:data <=32'hFFEFFFB9;
14'd5466:data <=32'hFFE0FFC2;14'd5467:data <=32'hFFD6FFCE;14'd5468:data <=32'hFFD1FFDC;
14'd5469:data <=32'hFFD1FFEA;14'd5470:data <=32'hFFD5FFF6;14'd5471:data <=32'hFFDBFFFF;
14'd5472:data <=32'hFFE40005;14'd5473:data <=32'hFFED0008;14'd5474:data <=32'hFFF50008;
14'd5475:data <=32'hFFFD0006;14'd5476:data <=32'h00030002;14'd5477:data <=32'h0008FFFB;
14'd5478:data <=32'h000BFFF4;14'd5479:data <=32'h000BFFEC;14'd5480:data <=32'h0009FFE3;
14'd5481:data <=32'h0003FFDB;14'd5482:data <=32'hFFFBFFD5;14'd5483:data <=32'hFFF1FFD1;
14'd5484:data <=32'hFFE6FFD0;14'd5485:data <=32'hFFDCFFD3;14'd5486:data <=32'hFFD3FFD7;
14'd5487:data <=32'hFFCCFFDE;14'd5488:data <=32'hFFC7FFE3;14'd5489:data <=32'hFFC2FFE9;
14'd5490:data <=32'hFFBDFFEF;14'd5491:data <=32'hFFB8FFF6;14'd5492:data <=32'hFFB1FFFE;
14'd5493:data <=32'hFFAC0009;14'd5494:data <=32'hFFA80017;14'd5495:data <=32'hFFA70027;
14'd5496:data <=32'hFFAB0039;14'd5497:data <=32'hFFB3004A;14'd5498:data <=32'hFFBF0058;
14'd5499:data <=32'hFFCF0064;14'd5500:data <=32'hFFE0006C;14'd5501:data <=32'hFFF20070;
14'd5502:data <=32'h00060071;14'd5503:data <=32'h0019006F;14'd5504:data <=32'hFFD9001A;
14'd5505:data <=32'hFFD70031;14'd5506:data <=32'hFFE4004A;14'd5507:data <=32'h002F0061;
14'd5508:data <=32'h00570048;14'd5509:data <=32'h005C0031;14'd5510:data <=32'h005A001A;
14'd5511:data <=32'h00520007;14'd5512:data <=32'h0046FFFA;14'd5513:data <=32'h0038FFF3;
14'd5514:data <=32'h002CFFF1;14'd5515:data <=32'h0023FFF3;14'd5516:data <=32'h001CFFF7;
14'd5517:data <=32'h0019FFFB;14'd5518:data <=32'h00180000;14'd5519:data <=32'h00190003;
14'd5520:data <=32'h001B0006;14'd5521:data <=32'h001F0007;14'd5522:data <=32'h00240007;
14'd5523:data <=32'h002B0005;14'd5524:data <=32'h0030FFFF;14'd5525:data <=32'h0035FFF7;
14'd5526:data <=32'h0036FFED;14'd5527:data <=32'h0034FFE1;14'd5528:data <=32'h002DFFD7;
14'd5529:data <=32'h0024FFD0;14'd5530:data <=32'h0019FFCC;14'd5531:data <=32'h000EFFCD;
14'd5532:data <=32'h0005FFD0;14'd5533:data <=32'hFFFFFFD4;14'd5534:data <=32'hFFFAFFD9;
14'd5535:data <=32'hFFF9FFDE;14'd5536:data <=32'hFFF7FFE1;14'd5537:data <=32'hFFF7FFE5;
14'd5538:data <=32'hFFF6FFE7;14'd5539:data <=32'hFFF5FFEA;14'd5540:data <=32'hFFF4FFED;
14'd5541:data <=32'hFFF5FFF1;14'd5542:data <=32'hFFF7FFF3;14'd5543:data <=32'hFFFAFFF6;
14'd5544:data <=32'hFFFEFFF6;14'd5545:data <=32'h0002FFF5;14'd5546:data <=32'h0005FFF2;
14'd5547:data <=32'h0008FFEF;14'd5548:data <=32'h0009FFEB;14'd5549:data <=32'h000AFFE6;
14'd5550:data <=32'h000AFFE1;14'd5551:data <=32'h0009FFDA;14'd5552:data <=32'h0007FFD2;
14'd5553:data <=32'h0002FFC9;14'd5554:data <=32'hFFFAFFBF;14'd5555:data <=32'hFFEDFFB7;
14'd5556:data <=32'hFFDCFFB1;14'd5557:data <=32'hFFC7FFB1;14'd5558:data <=32'hFFB2FFB7;
14'd5559:data <=32'hFF9DFFC4;14'd5560:data <=32'hFF8CFFD7;14'd5561:data <=32'hFF81FFEF;
14'd5562:data <=32'hFF7C0009;14'd5563:data <=32'hFF7D0024;14'd5564:data <=32'hFF85003D;
14'd5565:data <=32'hFF920054;14'd5566:data <=32'hFFA40068;14'd5567:data <=32'hFFB90077;
14'd5568:data <=32'hFFCB002A;14'd5569:data <=32'hFFC9003A;14'd5570:data <=32'hFFC6004F;
14'd5571:data <=32'hFFCD0079;14'd5572:data <=32'hFFFF0073;14'd5573:data <=32'h00120069;
14'd5574:data <=32'h0020005D;14'd5575:data <=32'h0029004E;14'd5576:data <=32'h002E0041;
14'd5577:data <=32'h002F0037;14'd5578:data <=32'h002F002F;14'd5579:data <=32'h002F0029;
14'd5580:data <=32'h00300024;14'd5581:data <=32'h0031001F;14'd5582:data <=32'h00330019;
14'd5583:data <=32'h00330012;14'd5584:data <=32'h0032000C;14'd5585:data <=32'h00300007;
14'd5586:data <=32'h002E0003;14'd5587:data <=32'h002B0000;14'd5588:data <=32'h002AFFFD;
14'd5589:data <=32'h0028FFF9;14'd5590:data <=32'h0026FFF6;14'd5591:data <=32'h0023FFF2;
14'd5592:data <=32'h001FFFEF;14'd5593:data <=32'h0019FFED;14'd5594:data <=32'h0014FFEE;
14'd5595:data <=32'h0010FFF1;14'd5596:data <=32'h000EFFF5;14'd5597:data <=32'h000FFFFA;
14'd5598:data <=32'h0012FFFD;14'd5599:data <=32'h0017FFFD;14'd5600:data <=32'h001CFFFA;
14'd5601:data <=32'h001FFFF5;14'd5602:data <=32'h0020FFEF;14'd5603:data <=32'h001EFFE8;
14'd5604:data <=32'h001AFFE3;14'd5605:data <=32'h0014FFE0;14'd5606:data <=32'h000FFFDF;
14'd5607:data <=32'h0009FFDF;14'd5608:data <=32'h0005FFE1;14'd5609:data <=32'h0002FFE4;
14'd5610:data <=32'h0000FFE7;14'd5611:data <=32'h0000FFEA;14'd5612:data <=32'h0001FFEE;
14'd5613:data <=32'h0004FFF0;14'd5614:data <=32'h0009FFF2;14'd5615:data <=32'h000EFFF1;
14'd5616:data <=32'h0015FFEE;14'd5617:data <=32'h001BFFE6;14'd5618:data <=32'h001EFFDB;
14'd5619:data <=32'h001DFFCD;14'd5620:data <=32'h0017FFBE;14'd5621:data <=32'h000BFFB1;
14'd5622:data <=32'hFFFAFFA7;14'd5623:data <=32'hFFE6FFA3;14'd5624:data <=32'hFFD1FFA4;
14'd5625:data <=32'hFFBDFFAC;14'd5626:data <=32'hFFACFFB9;14'd5627:data <=32'hFF9EFFC8;
14'd5628:data <=32'hFF95FFDA;14'd5629:data <=32'hFF8EFFED;14'd5630:data <=32'hFF8C0000;
14'd5631:data <=32'hFF8E0014;14'd5632:data <=32'hFF8E0005;14'd5633:data <=32'hFF86001E;
14'd5634:data <=32'hFF85002F;14'd5635:data <=32'hFF92001D;14'd5636:data <=32'hFFB20025;
14'd5637:data <=32'hFFB9002D;14'd5638:data <=32'hFFBF0033;14'd5639:data <=32'hFFC40038;
14'd5640:data <=32'hFFC8003F;14'd5641:data <=32'hFFCE0047;14'd5642:data <=32'hFFD5004F;
14'd5643:data <=32'hFFDF0059;14'd5644:data <=32'hFFEE0060;14'd5645:data <=32'hFFFF0063;
14'd5646:data <=32'h00110063;14'd5647:data <=32'h0023005D;14'd5648:data <=32'h00320052;
14'd5649:data <=32'h003E0044;14'd5650:data <=32'h00450035;14'd5651:data <=32'h00490025;
14'd5652:data <=32'h004A0016;14'd5653:data <=32'h00470007;14'd5654:data <=32'h0041FFFA;
14'd5655:data <=32'h0039FFEE;14'd5656:data <=32'h002EFFE6;14'd5657:data <=32'h0020FFE1;
14'd5658:data <=32'h0012FFE1;14'd5659:data <=32'h0005FFE6;14'd5660:data <=32'hFFFCFFEF;
14'd5661:data <=32'hFFF7FFFA;14'd5662:data <=32'hFFF70006;14'd5663:data <=32'hFFFC0010;
14'd5664:data <=32'h00040017;14'd5665:data <=32'h000D001A;14'd5666:data <=32'h00170019;
14'd5667:data <=32'h001E0015;14'd5668:data <=32'h00240010;14'd5669:data <=32'h0028000A;
14'd5670:data <=32'h002A0004;14'd5671:data <=32'h002AFFFF;14'd5672:data <=32'h002AFFFA;
14'd5673:data <=32'h002AFFF5;14'd5674:data <=32'h0029FFF0;14'd5675:data <=32'h0027FFEB;
14'd5676:data <=32'h0024FFE8;14'd5677:data <=32'h0022FFE5;14'd5678:data <=32'h0020FFE3;
14'd5679:data <=32'h001EFFE2;14'd5680:data <=32'h001EFFE0;14'd5681:data <=32'h001FFFDD;
14'd5682:data <=32'h001FFFD8;14'd5683:data <=32'h001EFFD1;14'd5684:data <=32'h001BFFC9;
14'd5685:data <=32'h0014FFC1;14'd5686:data <=32'h000BFFBA;14'd5687:data <=32'hFFFFFFB6;
14'd5688:data <=32'hFFF2FFB7;14'd5689:data <=32'hFFE7FFBA;14'd5690:data <=32'hFFDEFFC0;
14'd5691:data <=32'hFFD7FFC7;14'd5692:data <=32'hFFD2FFCE;14'd5693:data <=32'hFFCFFFD4;
14'd5694:data <=32'hFFCCFFD8;14'd5695:data <=32'hFFC9FFDD;14'd5696:data <=32'hFFA7FFA7;
14'd5697:data <=32'hFF8DFFB6;14'd5698:data <=32'hFF83FFCD;14'd5699:data <=32'hFFC1FFDE;
14'd5700:data <=32'hFFD8FFDC;14'd5701:data <=32'hFFD1FFDB;14'd5702:data <=32'hFFC8FFDB;
14'd5703:data <=32'hFFBDFFDD;14'd5704:data <=32'hFFB0FFE4;14'd5705:data <=32'hFFA4FFF0;
14'd5706:data <=32'hFF9A0001;14'd5707:data <=32'hFF960016;14'd5708:data <=32'hFF98002D;
14'd5709:data <=32'hFFA20044;14'd5710:data <=32'hFFB10056;14'd5711:data <=32'hFFC50063;
14'd5712:data <=32'hFFDB006B;14'd5713:data <=32'hFFF1006C;14'd5714:data <=32'h00070069;
14'd5715:data <=32'h00190061;14'd5716:data <=32'h00290056;14'd5717:data <=32'h00360048;
14'd5718:data <=32'h003E0037;14'd5719:data <=32'h00430026;14'd5720:data <=32'h00430014;
14'd5721:data <=32'h003D0003;14'd5722:data <=32'h0033FFF6;14'd5723:data <=32'h0026FFEE;
14'd5724:data <=32'h0018FFEA;14'd5725:data <=32'h000CFFEC;14'd5726:data <=32'h0002FFF1;
14'd5727:data <=32'hFFFBFFF8;14'd5728:data <=32'hFFF80000;14'd5729:data <=32'hFFF70007;
14'd5730:data <=32'hFFF8000D;14'd5731:data <=32'hFFFA0012;14'd5732:data <=32'hFFFB0017;
14'd5733:data <=32'hFFFE001C;14'd5734:data <=32'h00020021;14'd5735:data <=32'h00070026;
14'd5736:data <=32'h000F002A;14'd5737:data <=32'h0018002D;14'd5738:data <=32'h0023002D;
14'd5739:data <=32'h002E0029;14'd5740:data <=32'h00380024;14'd5741:data <=32'h0041001C;
14'd5742:data <=32'h00490012;14'd5743:data <=32'h004E0006;14'd5744:data <=32'h0052FFFA;
14'd5745:data <=32'h0053FFEC;14'd5746:data <=32'h0052FFDE;14'd5747:data <=32'h004EFFCE;
14'd5748:data <=32'h0046FFBF;14'd5749:data <=32'h003AFFB2;14'd5750:data <=32'h002AFFA8;
14'd5751:data <=32'h0017FFA3;14'd5752:data <=32'h0004FFA4;14'd5753:data <=32'hFFF3FFAA;
14'd5754:data <=32'hFFE6FFB5;14'd5755:data <=32'hFFDDFFC1;14'd5756:data <=32'hFFDAFFCE;
14'd5757:data <=32'hFFDBFFD9;14'd5758:data <=32'hFFDEFFE1;14'd5759:data <=32'hFFE3FFE5;
14'd5760:data <=32'hFFFFFFA5;14'd5761:data <=32'hFFEBFF9E;14'd5762:data <=32'hFFD5FFA6;
14'd5763:data <=32'hFFD8FFDE;14'd5764:data <=32'hFFF4FFDC;14'd5765:data <=32'hFFF3FFD6;
14'd5766:data <=32'hFFEFFFD0;14'd5767:data <=32'hFFE8FFCA;14'd5768:data <=32'hFFDDFFC6;
14'd5769:data <=32'hFFCFFFC6;14'd5770:data <=32'hFFBFFFCC;14'd5771:data <=32'hFFB2FFD6;
14'd5772:data <=32'hFFA7FFE6;14'd5773:data <=32'hFFA2FFF8;14'd5774:data <=32'hFFA3000A;
14'd5775:data <=32'hFFA8001A;14'd5776:data <=32'hFFB10029;14'd5777:data <=32'hFFBB0033;
14'd5778:data <=32'hFFC7003B;14'd5779:data <=32'hFFD20040;14'd5780:data <=32'hFFDE0044;
14'd5781:data <=32'hFFEA0045;14'd5782:data <=32'hFFF60044;14'd5783:data <=32'h00010040;
14'd5784:data <=32'h000B003A;14'd5785:data <=32'h00130032;14'd5786:data <=32'h00170029;
14'd5787:data <=32'h00190021;14'd5788:data <=32'h00180019;14'd5789:data <=32'h00170014;
14'd5790:data <=32'h0015000F;14'd5791:data <=32'h0013000C;14'd5792:data <=32'h00110008;
14'd5793:data <=32'h000F0005;14'd5794:data <=32'h000C0001;14'd5795:data <=32'h0007FFFD;
14'd5796:data <=32'hFFFFFFFB;14'd5797:data <=32'hFFF6FFFC;14'd5798:data <=32'hFFED0001;
14'd5799:data <=32'hFFE7000A;14'd5800:data <=32'hFFE20016;14'd5801:data <=32'hFFE20023;
14'd5802:data <=32'hFFE70031;14'd5803:data <=32'hFFF0003D;14'd5804:data <=32'hFFFD0046;
14'd5805:data <=32'h000C004C;14'd5806:data <=32'h001D004F;14'd5807:data <=32'h002F004D;
14'd5808:data <=32'h00400047;14'd5809:data <=32'h0051003D;14'd5810:data <=32'h005F002E;
14'd5811:data <=32'h006A001C;14'd5812:data <=32'h00710006;14'd5813:data <=32'h0072FFEF;
14'd5814:data <=32'h006BFFD8;14'd5815:data <=32'h005FFFC4;14'd5816:data <=32'h004EFFB5;
14'd5817:data <=32'h003BFFAC;14'd5818:data <=32'h0028FFAA;14'd5819:data <=32'h0017FFAC;
14'd5820:data <=32'h000BFFB2;14'd5821:data <=32'h0002FFB9;14'd5822:data <=32'hFFFCFFBF;
14'd5823:data <=32'hFFF8FFC5;14'd5824:data <=32'h000CFFD1;14'd5825:data <=32'h000AFFCB;
14'd5826:data <=32'h0000FFC2;14'd5827:data <=32'hFFE9FFB4;14'd5828:data <=32'hFFFCFFB8;
14'd5829:data <=32'hFFF5FFB8;14'd5830:data <=32'hFFEEFFB9;14'd5831:data <=32'hFFE6FFBB;
14'd5832:data <=32'hFFDDFFBD;14'd5833:data <=32'hFFD3FFC1;14'd5834:data <=32'hFFC9FFC8;
14'd5835:data <=32'hFFC0FFD1;14'd5836:data <=32'hFFBBFFDE;14'd5837:data <=32'hFFBAFFEC;
14'd5838:data <=32'hFFBCFFF9;14'd5839:data <=32'hFFC20004;14'd5840:data <=32'hFFCA000B;
14'd5841:data <=32'hFFD3000E;14'd5842:data <=32'hFFD9000F;14'd5843:data <=32'hFFDE000E;
14'd5844:data <=32'hFFE0000C;14'd5845:data <=32'hFFE0000C;14'd5846:data <=32'hFFE0000D;
14'd5847:data <=32'hFFE1000E;14'd5848:data <=32'hFFE10010;14'd5849:data <=32'hFFE10012;
14'd5850:data <=32'hFFE20014;14'd5851:data <=32'hFFE20017;14'd5852:data <=32'hFFE4001A;
14'd5853:data <=32'hFFE6001F;14'd5854:data <=32'hFFEB0023;14'd5855:data <=32'hFFF10026;
14'd5856:data <=32'hFFF80027;14'd5857:data <=32'h00010025;14'd5858:data <=32'h00080020;
14'd5859:data <=32'h000D0018;14'd5860:data <=32'h000E000E;14'd5861:data <=32'h000A0006;
14'd5862:data <=32'h0003FFFF;14'd5863:data <=32'hFFFAFFFC;14'd5864:data <=32'hFFF0FFFE;
14'd5865:data <=32'hFFE60003;14'd5866:data <=32'hFFE0000B;14'd5867:data <=32'hFFDC0016;
14'd5868:data <=32'hFFDC0022;14'd5869:data <=32'hFFDF002D;14'd5870:data <=32'hFFE50038;
14'd5871:data <=32'hFFED0041;14'd5872:data <=32'hFFF80049;14'd5873:data <=32'h0005004F;
14'd5874:data <=32'h00140052;14'd5875:data <=32'h00250051;14'd5876:data <=32'h0035004C;
14'd5877:data <=32'h00430042;14'd5878:data <=32'h004E0035;14'd5879:data <=32'h00550027;
14'd5880:data <=32'h00580018;14'd5881:data <=32'h0058000C;14'd5882:data <=32'h00560001;
14'd5883:data <=32'h0054FFF8;14'd5884:data <=32'h0053FFF0;14'd5885:data <=32'h0053FFE8;
14'd5886:data <=32'h0052FFDE;14'd5887:data <=32'h0050FFD3;14'd5888:data <=32'h0016FFCA;
14'd5889:data <=32'h0013FFCB;14'd5890:data <=32'h0017FFCA;14'd5891:data <=32'h0046FFB3;
14'd5892:data <=32'h0054FFA6;14'd5893:data <=32'h0042FF98;14'd5894:data <=32'h002FFF8E;
14'd5895:data <=32'h0019FF89;14'd5896:data <=32'h0003FF88;14'd5897:data <=32'hFFEDFF8B;
14'd5898:data <=32'hFFD7FF94;14'd5899:data <=32'hFFC4FFA2;14'd5900:data <=32'hFFB6FFB5;
14'd5901:data <=32'hFFAEFFCB;14'd5902:data <=32'hFFADFFE1;14'd5903:data <=32'hFFB3FFF5;
14'd5904:data <=32'hFFBE0004;14'd5905:data <=32'hFFCB000E;14'd5906:data <=32'hFFD90012;
14'd5907:data <=32'hFFE50011;14'd5908:data <=32'hFFEE000D;14'd5909:data <=32'hFFF40008;
14'd5910:data <=32'hFFF70002;14'd5911:data <=32'hFFF8FFFC;14'd5912:data <=32'hFFF6FFF7;
14'd5913:data <=32'hFFF4FFF3;14'd5914:data <=32'hFFEFFFEF;14'd5915:data <=32'hFFEAFFEE;
14'd5916:data <=32'hFFE3FFEF;14'd5917:data <=32'hFFDDFFF3;14'd5918:data <=32'hFFD8FFF8;
14'd5919:data <=32'hFFD60000;14'd5920:data <=32'hFFD70009;14'd5921:data <=32'hFFDA000F;
14'd5922:data <=32'hFFE00013;14'd5923:data <=32'hFFE60015;14'd5924:data <=32'hFFEA0015;
14'd5925:data <=32'hFFED0012;14'd5926:data <=32'hFFEE000F;14'd5927:data <=32'hFFED000D;
14'd5928:data <=32'hFFEA000D;14'd5929:data <=32'hFFE8000F;14'd5930:data <=32'hFFE60012;
14'd5931:data <=32'hFFE60016;14'd5932:data <=32'hFFE70019;14'd5933:data <=32'hFFE9001C;
14'd5934:data <=32'hFFEB001F;14'd5935:data <=32'hFFEC0021;14'd5936:data <=32'hFFED0023;
14'd5937:data <=32'hFFEF0026;14'd5938:data <=32'hFFF00029;14'd5939:data <=32'hFFF3002D;
14'd5940:data <=32'hFFF70031;14'd5941:data <=32'hFFFB0033;14'd5942:data <=32'hFFFF0036;
14'd5943:data <=32'h00030038;14'd5944:data <=32'h0007003B;14'd5945:data <=32'h000C003F;
14'd5946:data <=32'h00120044;14'd5947:data <=32'h001C004A;14'd5948:data <=32'h002A004E;
14'd5949:data <=32'h003B004E;14'd5950:data <=32'h004F004A;14'd5951:data <=32'h0062003F;
14'd5952:data <=32'h0046FFF5;14'd5953:data <=32'h0048FFF0;14'd5954:data <=32'h0048FFF3;
14'd5955:data <=32'h006B001A;14'd5956:data <=32'h008B0004;14'd5957:data <=32'h008AFFE9;
14'd5958:data <=32'h0083FFD0;14'd5959:data <=32'h0076FFB8;14'd5960:data <=32'h0065FFA4;
14'd5961:data <=32'h004FFF94;14'd5962:data <=32'h0036FF89;14'd5963:data <=32'h001CFF86;
14'd5964:data <=32'h0001FF89;14'd5965:data <=32'hFFEAFF94;14'd5966:data <=32'hFFD9FFA4;
14'd5967:data <=32'hFFCEFFB6;14'd5968:data <=32'hFFC9FFC8;14'd5969:data <=32'hFFCAFFD8;
14'd5970:data <=32'hFFCEFFE5;14'd5971:data <=32'hFFD3FFEE;14'd5972:data <=32'hFFD9FFF4;
14'd5973:data <=32'hFFDEFFF9;14'd5974:data <=32'hFFE3FFFC;14'd5975:data <=32'hFFE8FFFF;
14'd5976:data <=32'hFFED0000;14'd5977:data <=32'hFFF2FFFF;14'd5978:data <=32'hFFF7FFFD;
14'd5979:data <=32'hFFFAFFFA;14'd5980:data <=32'hFFFBFFF6;14'd5981:data <=32'hFFFAFFF2;
14'd5982:data <=32'hFFF8FFEF;14'd5983:data <=32'hFFF6FFED;14'd5984:data <=32'hFFF3FFEC;
14'd5985:data <=32'hFFF1FFEC;14'd5986:data <=32'hFFEFFFEB;14'd5987:data <=32'hFFECFFEA;
14'd5988:data <=32'hFFE9FFE8;14'd5989:data <=32'hFFE3FFE7;14'd5990:data <=32'hFFDDFFE7;
14'd5991:data <=32'hFFD5FFEA;14'd5992:data <=32'hFFCDFFF0;14'd5993:data <=32'hFFC7FFF8;
14'd5994:data <=32'hFFC40003;14'd5995:data <=32'hFFC5000F;14'd5996:data <=32'hFFC9001A;
14'd5997:data <=32'hFFD10022;14'd5998:data <=32'hFFD90027;14'd5999:data <=32'hFFE2002A;
14'd6000:data <=32'hFFE90029;14'd6001:data <=32'hFFF00026;14'd6002:data <=32'hFFF30023;
14'd6003:data <=32'hFFF60020;14'd6004:data <=32'hFFF6001C;14'd6005:data <=32'hFFF50019;
14'd6006:data <=32'hFFF30017;14'd6007:data <=32'hFFEE0016;14'd6008:data <=32'hFFE80018;
14'd6009:data <=32'hFFE2001F;14'd6010:data <=32'hFFDD0029;14'd6011:data <=32'hFFDC0037;
14'd6012:data <=32'hFFE00046;14'd6013:data <=32'hFFEA0056;14'd6014:data <=32'hFFFB0063;
14'd6015:data <=32'h0011006A;14'd6016:data <=32'h001B0049;14'd6017:data <=32'h002B004E;
14'd6018:data <=32'h0033004D;14'd6019:data <=32'h00260050;14'd6020:data <=32'h004F0049;
14'd6021:data <=32'h005A003B;14'd6022:data <=32'h0062002B;14'd6023:data <=32'h0067001A;
14'd6024:data <=32'h00690009;14'd6025:data <=32'h0067FFF7;14'd6026:data <=32'h0061FFE6;
14'd6027:data <=32'h0058FFD8;14'd6028:data <=32'h004CFFCD;14'd6029:data <=32'h003FFFC5;
14'd6030:data <=32'h0032FFC2;14'd6031:data <=32'h0027FFC2;14'd6032:data <=32'h001FFFC3;
14'd6033:data <=32'h0018FFC3;14'd6034:data <=32'h0013FFC3;14'd6035:data <=32'h000CFFC2;
14'd6036:data <=32'h0004FFC1;14'd6037:data <=32'hFFFBFFC3;14'd6038:data <=32'hFFF1FFC6;
14'd6039:data <=32'hFFE8FFCC;14'd6040:data <=32'hFFE1FFD4;14'd6041:data <=32'hFFDEFFDE;
14'd6042:data <=32'hFFDDFFE8;14'd6043:data <=32'hFFDFFFF1;14'd6044:data <=32'hFFE3FFF9;
14'd6045:data <=32'hFFE9FFFF;14'd6046:data <=32'hFFF00002;14'd6047:data <=32'hFFF70004;
14'd6048:data <=32'hFFFE0004;14'd6049:data <=32'h00050002;14'd6050:data <=32'h000CFFFC;
14'd6051:data <=32'h0011FFF4;14'd6052:data <=32'h0013FFE9;14'd6053:data <=32'h0012FFDE;
14'd6054:data <=32'h000BFFD3;14'd6055:data <=32'h0000FFCA;14'd6056:data <=32'hFFF3FFC5;
14'd6057:data <=32'hFFE4FFC5;14'd6058:data <=32'hFFD5FFCA;14'd6059:data <=32'hFFC9FFD3;
14'd6060:data <=32'hFFC1FFDF;14'd6061:data <=32'hFFBDFFEB;14'd6062:data <=32'hFFBDFFF7;
14'd6063:data <=32'hFFBF0001;14'd6064:data <=32'hFFC30009;14'd6065:data <=32'hFFC70010;
14'd6066:data <=32'hFFCB0015;14'd6067:data <=32'hFFCF0019;14'd6068:data <=32'hFFD4001C;
14'd6069:data <=32'hFFD8001D;14'd6070:data <=32'hFFDB001E;14'd6071:data <=32'hFFDD001E;
14'd6072:data <=32'hFFDD001E;14'd6073:data <=32'hFFDC001F;14'd6074:data <=32'hFFD80023;
14'd6075:data <=32'hFFD7002A;14'd6076:data <=32'hFFD60034;14'd6077:data <=32'hFFDA003F;
14'd6078:data <=32'hFFE2004A;14'd6079:data <=32'hFFEE0053;14'd6080:data <=32'hFFC20036;
14'd6081:data <=32'hFFC8004F;14'd6082:data <=32'hFFD8005D;14'd6083:data <=32'h00070040;
14'd6084:data <=32'h0028003E;14'd6085:data <=32'h002C0034;14'd6086:data <=32'h002D002C;
14'd6087:data <=32'h002D0026;14'd6088:data <=32'h002D0021;14'd6089:data <=32'h002D001D;
14'd6090:data <=32'h002D0019;14'd6091:data <=32'h002C0015;14'd6092:data <=32'h002C0014;
14'd6093:data <=32'h002C0013;14'd6094:data <=32'h002E0013;14'd6095:data <=32'h00320012;
14'd6096:data <=32'h00380010;14'd6097:data <=32'h003F000B;14'd6098:data <=32'h00460002;
14'd6099:data <=32'h004BFFF5;14'd6100:data <=32'h004AFFE6;14'd6101:data <=32'h0045FFD7;
14'd6102:data <=32'h003BFFC9;14'd6103:data <=32'h002DFFC0;14'd6104:data <=32'h001EFFBB;
14'd6105:data <=32'h000EFFBB;14'd6106:data <=32'h0000FFBF;14'd6107:data <=32'hFFF5FFC6;
14'd6108:data <=32'hFFECFFCF;14'd6109:data <=32'hFFE6FFD9;14'd6110:data <=32'hFFE3FFE4;
14'd6111:data <=32'hFFE3FFEF;14'd6112:data <=32'hFFE6FFF9;14'd6113:data <=32'hFFED0002;
14'd6114:data <=32'hFFF60008;14'd6115:data <=32'h0001000B;14'd6116:data <=32'h000C0009;
14'd6117:data <=32'h00160002;14'd6118:data <=32'h001DFFF9;14'd6119:data <=32'h0020FFEE;
14'd6120:data <=32'h001FFFE2;14'd6121:data <=32'h001AFFD8;14'd6122:data <=32'h0013FFD0;
14'd6123:data <=32'h000AFFCB;14'd6124:data <=32'h0002FFC8;14'd6125:data <=32'hFFFAFFC7;
14'd6126:data <=32'hFFF3FFC6;14'd6127:data <=32'hFFECFFC5;14'd6128:data <=32'hFFE3FFC5;
14'd6129:data <=32'hFFDBFFC5;14'd6130:data <=32'hFFD0FFC7;14'd6131:data <=32'hFFC6FFCC;
14'd6132:data <=32'hFFBCFFD3;14'd6133:data <=32'hFFB3FFDC;14'd6134:data <=32'hFFABFFE7;
14'd6135:data <=32'hFFA6FFF3;14'd6136:data <=32'hFFA30001;14'd6137:data <=32'hFFA2000E;
14'd6138:data <=32'hFFA2001D;14'd6139:data <=32'hFFA5002C;14'd6140:data <=32'hFFAB003C;
14'd6141:data <=32'hFFB5004C;14'd6142:data <=32'hFFC40059;14'd6143:data <=32'hFFD60062;
14'd6144:data <=32'hFFBFFFFD;14'd6145:data <=32'hFFB30011;14'd6146:data <=32'hFFB2002C;
14'd6147:data <=32'hFFF2005A;14'd6148:data <=32'h001A0055;14'd6149:data <=32'h00240046;
14'd6150:data <=32'h00280037;14'd6151:data <=32'h0027002A;14'd6152:data <=32'h00240020;
14'd6153:data <=32'h00200019;14'd6154:data <=32'h001A0014;14'd6155:data <=32'h00150012;
14'd6156:data <=32'h000F0012;14'd6157:data <=32'h000A0015;14'd6158:data <=32'h0007001B;
14'd6159:data <=32'h00090022;14'd6160:data <=32'h000E002A;14'd6161:data <=32'h0017002F;
14'd6162:data <=32'h00230030;14'd6163:data <=32'h0030002C;14'd6164:data <=32'h003C0024;
14'd6165:data <=32'h00430018;14'd6166:data <=32'h00460009;14'd6167:data <=32'h0045FFFC;
14'd6168:data <=32'h0040FFF0;14'd6169:data <=32'h0039FFE7;14'd6170:data <=32'h0031FFE0;
14'd6171:data <=32'h0029FFDB;14'd6172:data <=32'h0021FFD9;14'd6173:data <=32'h0019FFD8;
14'd6174:data <=32'h0011FFD8;14'd6175:data <=32'h0009FFDA;14'd6176:data <=32'h0002FFDE;
14'd6177:data <=32'hFFFDFFE4;14'd6178:data <=32'hFFFBFFEB;14'd6179:data <=32'hFFFBFFF1;
14'd6180:data <=32'hFFFDFFF7;14'd6181:data <=32'h0001FFFB;14'd6182:data <=32'h0006FFFD;
14'd6183:data <=32'h000AFFFD;14'd6184:data <=32'h000DFFFC;14'd6185:data <=32'h0010FFFB;
14'd6186:data <=32'h0013FFFA;14'd6187:data <=32'h0017FFF9;14'd6188:data <=32'h001CFFF7;
14'd6189:data <=32'h0021FFF3;14'd6190:data <=32'h0027FFEC;14'd6191:data <=32'h002CFFE2;
14'd6192:data <=32'h002EFFD5;14'd6193:data <=32'h002BFFC5;14'd6194:data <=32'h0024FFB6;
14'd6195:data <=32'h0018FFA8;14'd6196:data <=32'h0006FF9D;14'd6197:data <=32'hFFF2FF97;
14'd6198:data <=32'hFFDDFF95;14'd6199:data <=32'hFFC7FF99;14'd6200:data <=32'hFFB2FFA1;
14'd6201:data <=32'hFF9EFFAE;14'd6202:data <=32'hFF8DFFC0;14'd6203:data <=32'hFF80FFD6;
14'd6204:data <=32'hFF78FFEF;14'd6205:data <=32'hFF76000B;14'd6206:data <=32'hFF7B0027;
14'd6207:data <=32'hFF880041;14'd6208:data <=32'hFFC0FFFD;14'd6209:data <=32'hFFB60008;
14'd6210:data <=32'hFFA80018;14'd6211:data <=32'hFF9F0047;14'd6212:data <=32'hFFCB0053;
14'd6213:data <=32'hFFDB0052;14'd6214:data <=32'hFFE8004F;14'd6215:data <=32'hFFF20049;
14'd6216:data <=32'hFFFA0045;14'd6217:data <=32'h00010040;14'd6218:data <=32'h0006003B;
14'd6219:data <=32'h000A0035;14'd6220:data <=32'h000D0030;14'd6221:data <=32'h000D002C;
14'd6222:data <=32'h000D0029;14'd6223:data <=32'h000D0028;14'd6224:data <=32'h000F0029;
14'd6225:data <=32'h0012002A;14'd6226:data <=32'h0017002A;14'd6227:data <=32'h001D0028;
14'd6228:data <=32'h00230023;14'd6229:data <=32'h0027001C;14'd6230:data <=32'h00280014;
14'd6231:data <=32'h0026000D;14'd6232:data <=32'h00220008;14'd6233:data <=32'h001F0006;
14'd6234:data <=32'h001B0006;14'd6235:data <=32'h001A0007;14'd6236:data <=32'h001A0007;
14'd6237:data <=32'h001B0008;14'd6238:data <=32'h001E0007;14'd6239:data <=32'h001F0004;
14'd6240:data <=32'h00200001;14'd6241:data <=32'h0020FFFE;14'd6242:data <=32'h001FFFFB;
14'd6243:data <=32'h001EFFF8;14'd6244:data <=32'h001DFFF6;14'd6245:data <=32'h001BFFF3;
14'd6246:data <=32'h0019FFF1;14'd6247:data <=32'h0015FFEF;14'd6248:data <=32'h0011FFEF;
14'd6249:data <=32'h000CFFEF;14'd6250:data <=32'h0009FFF4;14'd6251:data <=32'h0007FFFA;
14'd6252:data <=32'h00080001;14'd6253:data <=32'h000E0007;14'd6254:data <=32'h0017000B;
14'd6255:data <=32'h0023000C;14'd6256:data <=32'h00300006;14'd6257:data <=32'h003BFFFD;
14'd6258:data <=32'h0042FFEE;14'd6259:data <=32'h0045FFDD;14'd6260:data <=32'h0043FFCA;
14'd6261:data <=32'h003CFFB9;14'd6262:data <=32'h0030FFA9;14'd6263:data <=32'h0021FF9C;
14'd6264:data <=32'h000FFF93;14'd6265:data <=32'hFFFAFF8D;14'd6266:data <=32'hFFE5FF8C;
14'd6267:data <=32'hFFCEFF90;14'd6268:data <=32'hFFB8FF9A;14'd6269:data <=32'hFFA5FFA9;
14'd6270:data <=32'hFF96FFBD;14'd6271:data <=32'hFF8DFFD3;14'd6272:data <=32'hFFA0FFCF;
14'd6273:data <=32'hFF93FFDE;14'd6274:data <=32'hFF8BFFE9;14'd6275:data <=32'hFF93FFDB;
14'd6276:data <=32'hFFABFFEE;14'd6277:data <=32'hFFAAFFF6;14'd6278:data <=32'hFFA8FFFF;
14'd6279:data <=32'hFFA60009;14'd6280:data <=32'hFFA60015;14'd6281:data <=32'hFFA80023;
14'd6282:data <=32'hFFAE0030;14'd6283:data <=32'hFFB7003D;14'd6284:data <=32'hFFC20047;
14'd6285:data <=32'hFFCF004E;14'd6286:data <=32'hFFDC0053;14'd6287:data <=32'hFFEA0056;
14'd6288:data <=32'hFFF80056;14'd6289:data <=32'h00070054;14'd6290:data <=32'h0015004F;
14'd6291:data <=32'h00230045;14'd6292:data <=32'h002D0039;14'd6293:data <=32'h0033002A;
14'd6294:data <=32'h00340019;14'd6295:data <=32'h0030000B;14'd6296:data <=32'h0027FFFF;
14'd6297:data <=32'h001CFFF8;14'd6298:data <=32'h0010FFF7;14'd6299:data <=32'h0006FFF9;
14'd6300:data <=32'hFFFFFFFF;14'd6301:data <=32'hFFFB0006;14'd6302:data <=32'hFFFA000E;
14'd6303:data <=32'hFFFC0014;14'd6304:data <=32'hFFFF0019;14'd6305:data <=32'h0004001D;
14'd6306:data <=32'h00090020;14'd6307:data <=32'h00100021;14'd6308:data <=32'h00160020;
14'd6309:data <=32'h001D001E;14'd6310:data <=32'h00220019;14'd6311:data <=32'h00260014;
14'd6312:data <=32'h0027000D;14'd6313:data <=32'h00270007;14'd6314:data <=32'h00240003;
14'd6315:data <=32'h00210001;14'd6316:data <=32'h001E0001;14'd6317:data <=32'h001D0003;
14'd6318:data <=32'h001F0006;14'd6319:data <=32'h00240008;14'd6320:data <=32'h002A0007;
14'd6321:data <=32'h00310003;14'd6322:data <=32'h0037FFFC;14'd6323:data <=32'h003AFFF3;
14'd6324:data <=32'h003CFFE9;14'd6325:data <=32'h0039FFDE;14'd6326:data <=32'h0035FFD5;
14'd6327:data <=32'h0030FFCD;14'd6328:data <=32'h002AFFC6;14'd6329:data <=32'h0023FFC0;
14'd6330:data <=32'h001BFFBA;14'd6331:data <=32'h0012FFB6;14'd6332:data <=32'h0008FFB3;
14'd6333:data <=32'hFFFDFFB2;14'd6334:data <=32'hFFF3FFB4;14'd6335:data <=32'hFFEAFFB7;
14'd6336:data <=32'hFFDBFF88;14'd6337:data <=32'hFFC2FF8B;14'd6338:data <=32'hFFB5FF99;
14'd6339:data <=32'hFFE8FFB5;14'd6340:data <=32'hFFFBFFB8;14'd6341:data <=32'hFFF0FFB0;
14'd6342:data <=32'hFFE1FFAB;14'd6343:data <=32'hFFD0FFAA;14'd6344:data <=32'hFFBBFFAF;
14'd6345:data <=32'hFFA9FFBA;14'd6346:data <=32'hFF9AFFCA;14'd6347:data <=32'hFF8FFFDF;
14'd6348:data <=32'hFF8BFFF4;14'd6349:data <=32'hFF8B000B;14'd6350:data <=32'hFF8F0020;
14'd6351:data <=32'hFF990034;14'd6352:data <=32'hFFA60046;14'd6353:data <=32'hFFB80054;
14'd6354:data <=32'hFFCC005E;14'd6355:data <=32'hFFE30062;14'd6356:data <=32'hFFFA0060;
14'd6357:data <=32'h000E0057;14'd6358:data <=32'h001E0049;14'd6359:data <=32'h00290038;
14'd6360:data <=32'h002C0026;14'd6361:data <=32'h002A0016;14'd6362:data <=32'h00240009;
14'd6363:data <=32'h001B0000;14'd6364:data <=32'h0012FFFB;14'd6365:data <=32'h000AFFFA;
14'd6366:data <=32'h0002FFFA;14'd6367:data <=32'hFFFCFFFC;14'd6368:data <=32'hFFF6FFFF;
14'd6369:data <=32'hFFF00004;14'd6370:data <=32'hFFED0009;14'd6371:data <=32'hFFEA0010;
14'd6372:data <=32'hFFEA0017;14'd6373:data <=32'hFFEC0020;14'd6374:data <=32'hFFF00026;
14'd6375:data <=32'hFFF6002C;14'd6376:data <=32'hFFFD0030;14'd6377:data <=32'h00040033;
14'd6378:data <=32'h000B0034;14'd6379:data <=32'h00120035;14'd6380:data <=32'h00190036;
14'd6381:data <=32'h00220036;14'd6382:data <=32'h002C0034;14'd6383:data <=32'h00370030;
14'd6384:data <=32'h00420029;14'd6385:data <=32'h004C001E;14'd6386:data <=32'h00530011;
14'd6387:data <=32'h00560001;14'd6388:data <=32'h0054FFF0;14'd6389:data <=32'h004DFFE2;
14'd6390:data <=32'h0044FFD6;14'd6391:data <=32'h0039FFCF;14'd6392:data <=32'h002DFFCB;
14'd6393:data <=32'h0023FFCA;14'd6394:data <=32'h001AFFCB;14'd6395:data <=32'h0013FFCF;
14'd6396:data <=32'h000DFFD2;14'd6397:data <=32'h000AFFD6;14'd6398:data <=32'h0009FFDB;
14'd6399:data <=32'h000AFFDE;14'd6400:data <=32'h0032FFAE;14'd6401:data <=32'h0026FFA0;
14'd6402:data <=32'h0013FF9F;14'd6403:data <=32'h0009FFD5;14'd6404:data <=32'h0026FFD8;
14'd6405:data <=32'h0026FFCA;14'd6406:data <=32'h0021FFBC;14'd6407:data <=32'h0017FFAE;
14'd6408:data <=32'h0007FFA5;14'd6409:data <=32'hFFF4FFA0;14'd6410:data <=32'hFFE1FFA1;
14'd6411:data <=32'hFFCFFFA8;14'd6412:data <=32'hFFC0FFB1;14'd6413:data <=32'hFFB3FFBE;
14'd6414:data <=32'hFFA9FFCD;14'd6415:data <=32'hFFA2FFDD;14'd6416:data <=32'hFF9FFFEF;
14'd6417:data <=32'hFF9F0001;14'd6418:data <=32'hFFA40012;14'd6419:data <=32'hFFAD0022;
14'd6420:data <=32'hFFBA002E;14'd6421:data <=32'hFFC90036;14'd6422:data <=32'hFFD80039;
14'd6423:data <=32'hFFE50038;14'd6424:data <=32'hFFF00033;14'd6425:data <=32'hFFF8002E;
14'd6426:data <=32'hFFFD0028;14'd6427:data <=32'h00010024;14'd6428:data <=32'h0004001F;
14'd6429:data <=32'h0007001B;14'd6430:data <=32'h000A0017;14'd6431:data <=32'h000C0011;
14'd6432:data <=32'h000C000A;14'd6433:data <=32'h000A0003;14'd6434:data <=32'h0005FFFC;
14'd6435:data <=32'hFFFEFFF7;14'd6436:data <=32'hFFF5FFF5;14'd6437:data <=32'hFFECFFF7;
14'd6438:data <=32'hFFE3FFFB;14'd6439:data <=32'hFFDB0002;14'd6440:data <=32'hFFD5000B;
14'd6441:data <=32'hFFD20015;14'd6442:data <=32'hFFD00021;14'd6443:data <=32'hFFD2002E;
14'd6444:data <=32'hFFD7003C;14'd6445:data <=32'hFFDF004A;14'd6446:data <=32'hFFEC0056;
14'd6447:data <=32'hFFFE005F;14'd6448:data <=32'h00120063;14'd6449:data <=32'h00280061;
14'd6450:data <=32'h003E0059;14'd6451:data <=32'h004F004A;14'd6452:data <=32'h005C0038;
14'd6453:data <=32'h00620023;14'd6454:data <=32'h0063000F;14'd6455:data <=32'h005FFFFD;
14'd6456:data <=32'h0057FFEF;14'd6457:data <=32'h004EFFE4;14'd6458:data <=32'h0043FFDC;
14'd6459:data <=32'h0039FFD7;14'd6460:data <=32'h0030FFD5;14'd6461:data <=32'h0027FFD5;
14'd6462:data <=32'h001FFFD7;14'd6463:data <=32'h001AFFDB;14'd6464:data <=32'h0029FFEB;
14'd6465:data <=32'h002DFFE8;14'd6466:data <=32'h002CFFDE;14'd6467:data <=32'h001AFFCC;
14'd6468:data <=32'h0031FFD4;14'd6469:data <=32'h002FFFCC;14'd6470:data <=32'h002AFFC3;
14'd6471:data <=32'h0022FFBA;14'd6472:data <=32'h0016FFB4;14'd6473:data <=32'h0008FFB1;
14'd6474:data <=32'hFFFBFFB2;14'd6475:data <=32'hFFEFFFB7;14'd6476:data <=32'hFFE6FFBE;
14'd6477:data <=32'hFFE0FFC6;14'd6478:data <=32'hFFDCFFCD;14'd6479:data <=32'hFFD9FFD3;
14'd6480:data <=32'hFFD7FFD9;14'd6481:data <=32'hFFD5FFDF;14'd6482:data <=32'hFFD4FFE5;
14'd6483:data <=32'hFFD4FFEB;14'd6484:data <=32'hFFD5FFF0;14'd6485:data <=32'hFFD7FFF4;
14'd6486:data <=32'hFFD9FFF7;14'd6487:data <=32'hFFDAFFF8;14'd6488:data <=32'hFFDAFFF8;
14'd6489:data <=32'hFFD8FFFA;14'd6490:data <=32'hFFD5FFFE;14'd6491:data <=32'hFFD30004;
14'd6492:data <=32'hFFD3000C;14'd6493:data <=32'hFFD60014;14'd6494:data <=32'hFFDC001B;
14'd6495:data <=32'hFFE5001F;14'd6496:data <=32'hFFEF0020;14'd6497:data <=32'hFFF9001E;
14'd6498:data <=32'h00000017;14'd6499:data <=32'h0004000F;14'd6500:data <=32'h00050006;
14'd6501:data <=32'h0002FFFE;14'd6502:data <=32'hFFFDFFF8;14'd6503:data <=32'hFFF6FFF3;
14'd6504:data <=32'hFFEDFFF0;14'd6505:data <=32'hFFE4FFF0;14'd6506:data <=32'hFFD9FFF3;
14'd6507:data <=32'hFFCFFFF9;14'd6508:data <=32'hFFC60003;14'd6509:data <=32'hFFC00011;
14'd6510:data <=32'hFFBE0021;14'd6511:data <=32'hFFC00032;14'd6512:data <=32'hFFC80042;
14'd6513:data <=32'hFFD50050;14'd6514:data <=32'hFFE50059;14'd6515:data <=32'hFFF7005E;
14'd6516:data <=32'h0008005D;14'd6517:data <=32'h00170059;14'd6518:data <=32'h00230053;
14'd6519:data <=32'h002D004B;14'd6520:data <=32'h00350044;14'd6521:data <=32'h003C003D;
14'd6522:data <=32'h00420035;14'd6523:data <=32'h0048002D;14'd6524:data <=32'h004E0024;
14'd6525:data <=32'h0052001A;14'd6526:data <=32'h00540010;14'd6527:data <=32'h00550005;
14'd6528:data <=32'h001FFFEB;14'd6529:data <=32'h001DFFF1;14'd6530:data <=32'h0025FFF6;
14'd6531:data <=32'h005CFFEE;14'd6532:data <=32'h0073FFE9;14'd6533:data <=32'h006EFFD4;
14'd6534:data <=32'h0064FFC0;14'd6535:data <=32'h0055FFAE;14'd6536:data <=32'h0041FFA1;
14'd6537:data <=32'h002AFF9A;14'd6538:data <=32'h0013FF9A;14'd6539:data <=32'hFFFEFFA1;
14'd6540:data <=32'hFFEEFFAD;14'd6541:data <=32'hFFE3FFBA;14'd6542:data <=32'hFFDDFFC9;
14'd6543:data <=32'hFFDBFFD6;14'd6544:data <=32'hFFDDFFE1;14'd6545:data <=32'hFFE1FFEB;
14'd6546:data <=32'hFFE6FFF2;14'd6547:data <=32'hFFECFFF6;14'd6548:data <=32'hFFF3FFF7;
14'd6549:data <=32'hFFF9FFF7;14'd6550:data <=32'hFFFFFFF3;14'd6551:data <=32'h0002FFEC;
14'd6552:data <=32'h0002FFE5;14'd6553:data <=32'hFFFEFFDE;14'd6554:data <=32'hFFF6FFD9;
14'd6555:data <=32'hFFEDFFD8;14'd6556:data <=32'hFFE3FFDB;14'd6557:data <=32'hFFDBFFE1;
14'd6558:data <=32'hFFD7FFEA;14'd6559:data <=32'hFFD6FFF3;14'd6560:data <=32'hFFD8FFFA;
14'd6561:data <=32'hFFDC0000;14'd6562:data <=32'hFFE10003;14'd6563:data <=32'hFFE50005;
14'd6564:data <=32'hFFE90004;14'd6565:data <=32'hFFEB0003;14'd6566:data <=32'hFFEC0002;
14'd6567:data <=32'hFFED0000;14'd6568:data <=32'hFFEDFFFE;14'd6569:data <=32'hFFECFFFC;
14'd6570:data <=32'hFFEAFFFA;14'd6571:data <=32'hFFE7FFF9;14'd6572:data <=32'hFFE2FFF8;
14'd6573:data <=32'hFFDDFFFA;14'd6574:data <=32'hFFD7FFFD;14'd6575:data <=32'hFFD30003;
14'd6576:data <=32'hFFD00009;14'd6577:data <=32'hFFD00011;14'd6578:data <=32'hFFD10017;
14'd6579:data <=32'hFFD3001D;14'd6580:data <=32'hFFD50021;14'd6581:data <=32'hFFD50025;
14'd6582:data <=32'hFFD5002A;14'd6583:data <=32'hFFD50031;14'd6584:data <=32'hFFD5003B;
14'd6585:data <=32'hFFD90046;14'd6586:data <=32'hFFE00053;14'd6587:data <=32'hFFEC005F;
14'd6588:data <=32'hFFFB0068;14'd6589:data <=32'h000E006E;14'd6590:data <=32'h0023006E;
14'd6591:data <=32'h0037006B;14'd6592:data <=32'h00320014;14'd6593:data <=32'h00310015;
14'd6594:data <=32'h00300020;14'd6595:data <=32'h004C0057;14'd6596:data <=32'h00760052;
14'd6597:data <=32'h00850039;14'd6598:data <=32'h008D001C;14'd6599:data <=32'h008EFFFE;
14'd6600:data <=32'h0086FFE1;14'd6601:data <=32'h0077FFC8;14'd6602:data <=32'h0062FFB6;
14'd6603:data <=32'h004AFFAB;14'd6604:data <=32'h0033FFA7;14'd6605:data <=32'h001FFFA9;
14'd6606:data <=32'h000FFFAF;14'd6607:data <=32'h0001FFB8;14'd6608:data <=32'hFFF8FFC1;
14'd6609:data <=32'hFFF1FFCB;14'd6610:data <=32'hFFEDFFD5;14'd6611:data <=32'hFFEBFFDF;
14'd6612:data <=32'hFFEDFFE8;14'd6613:data <=32'hFFF0FFEF;14'd6614:data <=32'hFFF6FFF4;
14'd6615:data <=32'hFFFCFFF6;14'd6616:data <=32'h0002FFF4;14'd6617:data <=32'h0005FFF1;
14'd6618:data <=32'h0007FFED;14'd6619:data <=32'h0005FFE9;14'd6620:data <=32'h0003FFE6;
14'd6621:data <=32'h0000FFE5;14'd6622:data <=32'hFFFDFFE6;14'd6623:data <=32'hFFFCFFE7;
14'd6624:data <=32'hFFFCFFE7;14'd6625:data <=32'hFFFDFFE6;14'd6626:data <=32'hFFFCFFE3;
14'd6627:data <=32'hFFFAFFE0;14'd6628:data <=32'hFFF7FFDD;14'd6629:data <=32'hFFF0FFDA;
14'd6630:data <=32'hFFEAFFDA;14'd6631:data <=32'hFFE3FFDD;14'd6632:data <=32'hFFDDFFE1;
14'd6633:data <=32'hFFD9FFE6;14'd6634:data <=32'hFFD6FFEC;14'd6635:data <=32'hFFD5FFF2;
14'd6636:data <=32'hFFD5FFF8;14'd6637:data <=32'hFFD6FFFD;14'd6638:data <=32'hFFD80001;
14'd6639:data <=32'hFFDA0005;14'd6640:data <=32'hFFDE0008;14'd6641:data <=32'hFFE2000A;
14'd6642:data <=32'hFFE60009;14'd6643:data <=32'hFFE90005;14'd6644:data <=32'hFFE90000;
14'd6645:data <=32'hFFE6FFFB;14'd6646:data <=32'hFFDFFFF6;14'd6647:data <=32'hFFD4FFF5;
14'd6648:data <=32'hFFC7FFF8;14'd6649:data <=32'hFFBB0002;14'd6650:data <=32'hFFB20010;
14'd6651:data <=32'hFFAC0023;14'd6652:data <=32'hFFAD0038;14'd6653:data <=32'hFFB4004C;
14'd6654:data <=32'hFFC1005F;14'd6655:data <=32'hFFD1006E;14'd6656:data <=32'hFFF00047;
14'd6657:data <=32'hFFF60054;14'd6658:data <=32'hFFF8005C;14'd6659:data <=32'hFFE90067;
14'd6660:data <=32'h00150077;14'd6661:data <=32'h002B0072;14'd6662:data <=32'h00400066;
14'd6663:data <=32'h00500057;14'd6664:data <=32'h005B0044;14'd6665:data <=32'h0061002F;
14'd6666:data <=32'h0061001C;14'd6667:data <=32'h005D000C;14'd6668:data <=32'h00570000;
14'd6669:data <=32'h0051FFF7;14'd6670:data <=32'h004BFFEF;14'd6671:data <=32'h0046FFE8;
14'd6672:data <=32'h0040FFE1;14'd6673:data <=32'h003AFFDB;14'd6674:data <=32'h0032FFD4;
14'd6675:data <=32'h002AFFD0;14'd6676:data <=32'h0020FFCE;14'd6677:data <=32'h0017FFCE;
14'd6678:data <=32'h000FFFD0;14'd6679:data <=32'h0008FFD3;14'd6680:data <=32'h0003FFD7;
14'd6681:data <=32'hFFFEFFDA;14'd6682:data <=32'hFFF9FFDF;14'd6683:data <=32'hFFF5FFE3;
14'd6684:data <=32'hFFF3FFEB;14'd6685:data <=32'hFFF2FFF2;14'd6686:data <=32'hFFF5FFFA;
14'd6687:data <=32'hFFFB0001;14'd6688:data <=32'h00030004;14'd6689:data <=32'h000D0005;
14'd6690:data <=32'h00170000;14'd6691:data <=32'h001EFFF8;14'd6692:data <=32'h0022FFED;
14'd6693:data <=32'h0022FFE1;14'd6694:data <=32'h001DFFD6;14'd6695:data <=32'h0015FFCD;
14'd6696:data <=32'h000BFFC7;14'd6697:data <=32'h0000FFC4;14'd6698:data <=32'hFFF6FFC4;
14'd6699:data <=32'hFFEBFFC6;14'd6700:data <=32'hFFE2FFCA;14'd6701:data <=32'hFFDBFFD0;
14'd6702:data <=32'hFFD5FFD7;14'd6703:data <=32'hFFD1FFE0;14'd6704:data <=32'hFFCFFFE8;
14'd6705:data <=32'hFFD0FFF1;14'd6706:data <=32'hFFD4FFF6;14'd6707:data <=32'hFFD8FFFA;
14'd6708:data <=32'hFFDDFFFB;14'd6709:data <=32'hFFE0FFF8;14'd6710:data <=32'hFFE0FFF3;
14'd6711:data <=32'hFFDBFFEF;14'd6712:data <=32'hFFD4FFED;14'd6713:data <=32'hFFCAFFEF;
14'd6714:data <=32'hFFC0FFF5;14'd6715:data <=32'hFFB8FFFF;14'd6716:data <=32'hFFB3000B;
14'd6717:data <=32'hFFB10019;14'd6718:data <=32'hFFB40028;14'd6719:data <=32'hFFB90035;
14'd6720:data <=32'hFFA5000D;14'd6721:data <=32'hFF9B0026;14'd6722:data <=32'hFF9E003A;
14'd6723:data <=32'hFFCB0033;14'd6724:data <=32'hFFE90047;14'd6725:data <=32'hFFF30047;
14'd6726:data <=32'hFFFC0045;14'd6727:data <=32'h00040042;14'd6728:data <=32'h000A003D;
14'd6729:data <=32'h000D0039;14'd6730:data <=32'h000F0035;14'd6731:data <=32'h000F0034;
14'd6732:data <=32'h00110036;14'd6733:data <=32'h00150039;14'd6734:data <=32'h001C003C;
14'd6735:data <=32'h0027003D;14'd6736:data <=32'h0033003A;14'd6737:data <=32'h003E0033;
14'd6738:data <=32'h00480028;14'd6739:data <=32'h004F001A;14'd6740:data <=32'h0051000B;
14'd6741:data <=32'h0050FFFC;14'd6742:data <=32'h004CFFEE;14'd6743:data <=32'h0045FFE2;
14'd6744:data <=32'h003CFFD8;14'd6745:data <=32'h0030FFD0;14'd6746:data <=32'h0023FFCB;
14'd6747:data <=32'h0014FFC9;14'd6748:data <=32'h0006FFCC;14'd6749:data <=32'hFFF9FFD3;
14'd6750:data <=32'hFFF0FFDE;14'd6751:data <=32'hFFECFFEC;14'd6752:data <=32'hFFECFFF9;
14'd6753:data <=32'hFFF20005;14'd6754:data <=32'hFFFC000E;14'd6755:data <=32'h00070011;
14'd6756:data <=32'h00130010;14'd6757:data <=32'h001D000C;14'd6758:data <=32'h00240005;
14'd6759:data <=32'h0029FFFD;14'd6760:data <=32'h002BFFF4;14'd6761:data <=32'h002CFFEB;
14'd6762:data <=32'h002AFFE2;14'd6763:data <=32'h0028FFDB;14'd6764:data <=32'h0024FFD3;
14'd6765:data <=32'h001FFFCB;14'd6766:data <=32'h0018FFC4;14'd6767:data <=32'h0010FFC0;
14'd6768:data <=32'h0006FFBC;14'd6769:data <=32'hFFFDFFBB;14'd6770:data <=32'hFFF4FFBB;
14'd6771:data <=32'hFFEBFFBC;14'd6772:data <=32'hFFE4FFBD;14'd6773:data <=32'hFFDCFFBE;
14'd6774:data <=32'hFFD3FFC0;14'd6775:data <=32'hFFC9FFC3;14'd6776:data <=32'hFFBDFFC8;
14'd6777:data <=32'hFFB2FFD1;14'd6778:data <=32'hFFA7FFDD;14'd6779:data <=32'hFFA0FFEE;
14'd6780:data <=32'hFF9E0000;14'd6781:data <=32'hFFA10011;14'd6782:data <=32'hFFA80021;
14'd6783:data <=32'hFFB3002D;14'd6784:data <=32'hFFC3FFCB;14'd6785:data <=32'hFFAAFFD5;
14'd6786:data <=32'hFF99FFED;14'd6787:data <=32'hFFC2002E;14'd6788:data <=32'hFFE4003E;
14'd6789:data <=32'hFFEF003A;14'd6790:data <=32'hFFF80033;14'd6791:data <=32'hFFFD002B;
14'd6792:data <=32'hFFFF0022;14'd6793:data <=32'hFFFD001A;14'd6794:data <=32'hFFF70015;
14'd6795:data <=32'hFFEF0013;14'd6796:data <=32'hFFE70017;14'd6797:data <=32'hFFE20020;
14'd6798:data <=32'hFFE2002C;14'd6799:data <=32'hFFE60038;14'd6800:data <=32'hFFEF0043;
14'd6801:data <=32'hFFFC0049;14'd6802:data <=32'h000A004C;14'd6803:data <=32'h0019004A;
14'd6804:data <=32'h00260044;14'd6805:data <=32'h0031003B;14'd6806:data <=32'h003A0032;
14'd6807:data <=32'h00400026;14'd6808:data <=32'h00440019;14'd6809:data <=32'h0045000C;
14'd6810:data <=32'h0043FFFE;14'd6811:data <=32'h003DFFF2;14'd6812:data <=32'h0034FFE8;
14'd6813:data <=32'h0028FFE2;14'd6814:data <=32'h001CFFE0;14'd6815:data <=32'h0011FFE1;
14'd6816:data <=32'h0008FFE7;14'd6817:data <=32'h0003FFEE;14'd6818:data <=32'h0001FFF5;
14'd6819:data <=32'h0001FFFB;14'd6820:data <=32'h00020000;14'd6821:data <=32'h00040003;
14'd6822:data <=32'h00070006;14'd6823:data <=32'h00090009;14'd6824:data <=32'h000C000C;
14'd6825:data <=32'h0010000F;14'd6826:data <=32'h00160012;14'd6827:data <=32'h001F0013;
14'd6828:data <=32'h00280012;14'd6829:data <=32'h0032000D;14'd6830:data <=32'h003C0005;
14'd6831:data <=32'h0043FFFA;14'd6832:data <=32'h0048FFEC;14'd6833:data <=32'h0049FFDD;
14'd6834:data <=32'h0048FFCE;14'd6835:data <=32'h0043FFBE;14'd6836:data <=32'h003BFFAE;
14'd6837:data <=32'h002FFF9F;14'd6838:data <=32'h001FFF92;14'd6839:data <=32'h000BFF88;
14'd6840:data <=32'hFFF3FF82;14'd6841:data <=32'hFFD9FF83;14'd6842:data <=32'hFFBEFF8C;
14'd6843:data <=32'hFFA7FF9C;14'd6844:data <=32'hFF95FFB1;14'd6845:data <=32'hFF8AFFCA;
14'd6846:data <=32'hFF86FFE5;14'd6847:data <=32'hFF8AFFFD;14'd6848:data <=32'hFFDBFFD0;
14'd6849:data <=32'hFFCAFFCE;14'd6850:data <=32'hFFB2FFD3;14'd6851:data <=32'hFF910001;
14'd6852:data <=32'hFFB0001F;14'd6853:data <=32'hFFBC0026;14'd6854:data <=32'hFFC8002A;
14'd6855:data <=32'hFFD3002C;14'd6856:data <=32'hFFDD002A;14'd6857:data <=32'hFFE40024;
14'd6858:data <=32'hFFE70020;14'd6859:data <=32'hFFE7001B;14'd6860:data <=32'hFFE4001A;
14'd6861:data <=32'hFFE1001C;14'd6862:data <=32'hFFDF0021;14'd6863:data <=32'hFFE00027;
14'd6864:data <=32'hFFE5002E;14'd6865:data <=32'hFFEB0033;14'd6866:data <=32'hFFF30036;
14'd6867:data <=32'hFFFB0035;14'd6868:data <=32'h00020033;14'd6869:data <=32'h00080030;
14'd6870:data <=32'h000C002D;14'd6871:data <=32'h000F002A;14'd6872:data <=32'h00130028;
14'd6873:data <=32'h00160024;14'd6874:data <=32'h00190021;14'd6875:data <=32'h001B001D;
14'd6876:data <=32'h001C0018;14'd6877:data <=32'h001C0014;14'd6878:data <=32'h001B0011;
14'd6879:data <=32'h0019000E;14'd6880:data <=32'h0019000E;14'd6881:data <=32'h0019000C;
14'd6882:data <=32'h001A000B;14'd6883:data <=32'h001C0009;14'd6884:data <=32'h001C0004;
14'd6885:data <=32'h001B0000;14'd6886:data <=32'h0016FFFC;14'd6887:data <=32'h0011FFF9;
14'd6888:data <=32'h000AFFFB;14'd6889:data <=32'h0004FFFF;14'd6890:data <=32'h00000006;
14'd6891:data <=32'hFFFF000F;14'd6892:data <=32'h00030019;14'd6893:data <=32'h000B0021;
14'd6894:data <=32'h00150027;14'd6895:data <=32'h00220029;14'd6896:data <=32'h00310028;
14'd6897:data <=32'h003F0022;14'd6898:data <=32'h004C0018;14'd6899:data <=32'h0057000B;
14'd6900:data <=32'h0060FFFB;14'd6901:data <=32'h0065FFE7;14'd6902:data <=32'h0065FFD0;
14'd6903:data <=32'h005FFFBA;14'd6904:data <=32'h0052FFA4;14'd6905:data <=32'h0040FF91;
14'd6906:data <=32'h0028FF84;14'd6907:data <=32'h000EFF7E;14'd6908:data <=32'hFFF4FF80;
14'd6909:data <=32'hFFDCFF88;14'd6910:data <=32'hFFC9FF95;14'd6911:data <=32'hFFBBFFA4;
14'd6912:data <=32'hFFD5FFAF;14'd6913:data <=32'hFFC7FFB1;14'd6914:data <=32'hFFBAFFAF;
14'd6915:data <=32'hFFB9FFA1;14'd6916:data <=32'hFFC3FFBC;14'd6917:data <=32'hFFBBFFC4;
14'd6918:data <=32'hFFB5FFCE;14'd6919:data <=32'hFFB0FFD9;14'd6920:data <=32'hFFADFFE4;
14'd6921:data <=32'hFFABFFEF;14'd6922:data <=32'hFFAAFFF9;14'd6923:data <=32'hFFAB0003;
14'd6924:data <=32'hFFAB000F;14'd6925:data <=32'hFFAE001B;14'd6926:data <=32'hFFB30029;
14'd6927:data <=32'hFFBC0035;14'd6928:data <=32'hFFC90040;14'd6929:data <=32'hFFD90046;
14'd6930:data <=32'hFFEA0047;14'd6931:data <=32'hFFFA0043;14'd6932:data <=32'h0006003A;
14'd6933:data <=32'h000E0030;14'd6934:data <=32'h00120025;14'd6935:data <=32'h0012001B;
14'd6936:data <=32'h000F0013;14'd6937:data <=32'h000B000D;14'd6938:data <=32'h00060009;
14'd6939:data <=32'h00010007;14'd6940:data <=32'hFFFC0007;14'd6941:data <=32'hFFF7000A;
14'd6942:data <=32'hFFF3000D;14'd6943:data <=32'hFFF00013;14'd6944:data <=32'hFFF0001A;
14'd6945:data <=32'hFFF30020;14'd6946:data <=32'hFFF90026;14'd6947:data <=32'h00000029;
14'd6948:data <=32'h00090029;14'd6949:data <=32'h00110026;14'd6950:data <=32'h00150020;
14'd6951:data <=32'h0018001A;14'd6952:data <=32'h00160014;14'd6953:data <=32'h00130010;
14'd6954:data <=32'h000F000F;14'd6955:data <=32'h000B0011;14'd6956:data <=32'h000A0015;
14'd6957:data <=32'h000B001A;14'd6958:data <=32'h000E001F;14'd6959:data <=32'h00130023;
14'd6960:data <=32'h001A0025;14'd6961:data <=32'h00210026;14'd6962:data <=32'h002A0024;
14'd6963:data <=32'h00320022;14'd6964:data <=32'h003B001D;14'd6965:data <=32'h00430016;
14'd6966:data <=32'h004B000C;14'd6967:data <=32'h00510000;14'd6968:data <=32'h0053FFF2;
14'd6969:data <=32'h0051FFE3;14'd6970:data <=32'h004CFFD6;14'd6971:data <=32'h0043FFCA;
14'd6972:data <=32'h003AFFC3;14'd6973:data <=32'h0030FFBE;14'd6974:data <=32'h0027FFBB;
14'd6975:data <=32'h0021FFB8;14'd6976:data <=32'h001DFF8F;14'd6977:data <=32'h000AFF85;
14'd6978:data <=32'hFFFDFF87;14'd6979:data <=32'h0023FFA8;14'd6980:data <=32'h002DFFAF;
14'd6981:data <=32'h0022FFA2;14'd6982:data <=32'h0012FF98;14'd6983:data <=32'h0000FF92;
14'd6984:data <=32'hFFEDFF91;14'd6985:data <=32'hFFD9FF93;14'd6986:data <=32'hFFC6FF99;
14'd6987:data <=32'hFFB2FFA3;14'd6988:data <=32'hFFA1FFB3;14'd6989:data <=32'hFF94FFC6;
14'd6990:data <=32'hFF8AFFDD;14'd6991:data <=32'hFF88FFF7;14'd6992:data <=32'hFF8D0011;
14'd6993:data <=32'hFF990028;14'd6994:data <=32'hFFAA0039;14'd6995:data <=32'hFFC00044;
14'd6996:data <=32'hFFD50048;14'd6997:data <=32'hFFE80045;14'd6998:data <=32'hFFF8003E;
14'd6999:data <=32'h00040035;14'd7000:data <=32'h000C002A;14'd7001:data <=32'h0010001F;
14'd7002:data <=32'h00110015;14'd7003:data <=32'h0010000B;14'd7004:data <=32'h000C0002;
14'd7005:data <=32'h0006FFFB;14'd7006:data <=32'hFFFEFFF7;14'd7007:data <=32'hFFF5FFF5;
14'd7008:data <=32'hFFECFFF7;14'd7009:data <=32'hFFE5FFFC;14'd7010:data <=32'hFFE00004;
14'd7011:data <=32'hFFDF000B;14'd7012:data <=32'hFFDF0013;14'd7013:data <=32'hFFE10019;
14'd7014:data <=32'hFFE4001D;14'd7015:data <=32'hFFE70020;14'd7016:data <=32'hFFE90024;
14'd7017:data <=32'hFFEA0028;14'd7018:data <=32'hFFEC002C;14'd7019:data <=32'hFFF00032;
14'd7020:data <=32'hFFF50038;14'd7021:data <=32'hFFFD003E;14'd7022:data <=32'h00080041;
14'd7023:data <=32'h00130041;14'd7024:data <=32'h001F003F;14'd7025:data <=32'h00290039;
14'd7026:data <=32'h00310032;14'd7027:data <=32'h00370029;14'd7028:data <=32'h003B0020;
14'd7029:data <=32'h003D0017;14'd7030:data <=32'h003E000F;14'd7031:data <=32'h003D0007;
14'd7032:data <=32'h003AFFFF;14'd7033:data <=32'h0036FFF8;14'd7034:data <=32'h0031FFF3;
14'd7035:data <=32'h002BFFF2;14'd7036:data <=32'h0025FFF3;14'd7037:data <=32'h0023FFF6;
14'd7038:data <=32'h0024FFFB;14'd7039:data <=32'h0029FFFF;14'd7040:data <=32'h005AFFD9;
14'd7041:data <=32'h005AFFC7;14'd7042:data <=32'h004EFFBD;14'd7043:data <=32'h0037FFEB;
14'd7044:data <=32'h004FFFF3;14'd7045:data <=32'h0053FFE2;14'd7046:data <=32'h0052FFD0;
14'd7047:data <=32'h004CFFBF;14'd7048:data <=32'h0041FFAF;14'd7049:data <=32'h0034FFA2;
14'd7050:data <=32'h0023FF96;14'd7051:data <=32'h000FFF8F;14'd7052:data <=32'hFFFAFF8C;
14'd7053:data <=32'hFFE3FF8F;14'd7054:data <=32'hFFCDFF98;14'd7055:data <=32'hFFBAFFA7;
14'd7056:data <=32'hFFADFFBA;14'd7057:data <=32'hFFA6FFCF;14'd7058:data <=32'hFFA5FFE4;
14'd7059:data <=32'hFFA9FFF7;14'd7060:data <=32'hFFB20005;14'd7061:data <=32'hFFBB0010;
14'd7062:data <=32'hFFC60017;14'd7063:data <=32'hFFCF001C;14'd7064:data <=32'hFFD7001E;
14'd7065:data <=32'hFFE00020;14'd7066:data <=32'hFFE80020;14'd7067:data <=32'hFFF1001F;
14'd7068:data <=32'hFFF9001C;14'd7069:data <=32'hFFFE0016;14'd7070:data <=32'h00030010;
14'd7071:data <=32'h00050008;14'd7072:data <=32'h00040001;14'd7073:data <=32'h0002FFFB;
14'd7074:data <=32'hFFFDFFF6;14'd7075:data <=32'hFFF9FFF2;14'd7076:data <=32'hFFF3FFF0;
14'd7077:data <=32'hFFEDFFEE;14'd7078:data <=32'hFFE6FFED;14'd7079:data <=32'hFFDDFFEE;
14'd7080:data <=32'hFFD3FFF1;14'd7081:data <=32'hFFC9FFF8;14'd7082:data <=32'hFFC00002;
14'd7083:data <=32'hFFBA0011;14'd7084:data <=32'hFFB70021;14'd7085:data <=32'hFFBB0034;
14'd7086:data <=32'hFFC40045;14'd7087:data <=32'hFFD20053;14'd7088:data <=32'hFFE4005C;
14'd7089:data <=32'hFFF70060;14'd7090:data <=32'h00090060;14'd7091:data <=32'h001A005A;
14'd7092:data <=32'h00280052;14'd7093:data <=32'h00340047;14'd7094:data <=32'h003D003B;
14'd7095:data <=32'h0042002E;14'd7096:data <=32'h00440020;14'd7097:data <=32'h00430013;
14'd7098:data <=32'h003D0008;14'd7099:data <=32'h00350000;14'd7100:data <=32'h002CFFFC;
14'd7101:data <=32'h0024FFFE;14'd7102:data <=32'h001F0002;14'd7103:data <=32'h001E0009;
14'd7104:data <=32'h002C0019;14'd7105:data <=32'h00380019;14'd7106:data <=32'h003F000F;
14'd7107:data <=32'h0032FFF8;14'd7108:data <=32'h00470005;14'd7109:data <=32'h004BFFFB;
14'd7110:data <=32'h004BFFEF;14'd7111:data <=32'h0048FFE3;14'd7112:data <=32'h0043FFD9;
14'd7113:data <=32'h003DFFD0;14'd7114:data <=32'h0036FFC9;14'd7115:data <=32'h002EFFC2;
14'd7116:data <=32'h0024FFBC;14'd7117:data <=32'h0018FFB8;14'd7118:data <=32'h000DFFB7;
14'd7119:data <=32'h0001FFB9;14'd7120:data <=32'hFFF7FFBF;14'd7121:data <=32'hFFF0FFC5;
14'd7122:data <=32'hFFECFFCC;14'd7123:data <=32'hFFEAFFD2;14'd7124:data <=32'hFFEAFFD6;
14'd7125:data <=32'hFFE9FFD8;14'd7126:data <=32'hFFE6FFD9;14'd7127:data <=32'hFFE2FFDA;
14'd7128:data <=32'hFFDDFFDC;14'd7129:data <=32'hFFD7FFE1;14'd7130:data <=32'hFFD3FFE9;
14'd7131:data <=32'hFFD1FFF1;14'd7132:data <=32'hFFD2FFFA;14'd7133:data <=32'hFFD60003;
14'd7134:data <=32'hFFDC0009;14'd7135:data <=32'hFFE2000D;14'd7136:data <=32'hFFEA000F;
14'd7137:data <=32'hFFF1000F;14'd7138:data <=32'hFFF8000D;14'd7139:data <=32'hFFFE0009;
14'd7140:data <=32'h00040003;14'd7141:data <=32'h0006FFFB;14'd7142:data <=32'h0007FFF1;
14'd7143:data <=32'h0003FFE6;14'd7144:data <=32'hFFFBFFDD;14'd7145:data <=32'hFFEFFFD6;
14'd7146:data <=32'hFFE0FFD4;14'd7147:data <=32'hFFD0FFD6;14'd7148:data <=32'hFFC0FFDF;
14'd7149:data <=32'hFFB5FFEC;14'd7150:data <=32'hFFADFFFD;14'd7151:data <=32'hFFAB000E;
14'd7152:data <=32'hFFAD0020;14'd7153:data <=32'hFFB4002F;14'd7154:data <=32'hFFBD003C;
14'd7155:data <=32'hFFC80045;14'd7156:data <=32'hFFD3004D;14'd7157:data <=32'hFFDF0052;
14'd7158:data <=32'hFFEC0056;14'd7159:data <=32'hFFF90056;14'd7160:data <=32'h00060055;
14'd7161:data <=32'h00110052;14'd7162:data <=32'h001A004C;14'd7163:data <=32'h00220045;
14'd7164:data <=32'h0026003F;14'd7165:data <=32'h002A003B;14'd7166:data <=32'h002E0037;
14'd7167:data <=32'h00320035;14'd7168:data <=32'h000C000B;14'd7169:data <=32'h000B0017;
14'd7170:data <=32'h00170021;14'd7171:data <=32'h004F0027;14'd7172:data <=32'h0068002B;
14'd7173:data <=32'h006D0015;14'd7174:data <=32'h006B0001;14'd7175:data <=32'h0065FFED;
14'd7176:data <=32'h005AFFDD;14'd7177:data <=32'h004CFFD1;14'd7178:data <=32'h003EFFCA;
14'd7179:data <=32'h0030FFC7;14'd7180:data <=32'h0023FFC6;14'd7181:data <=32'h0017FFC7;
14'd7182:data <=32'h000DFFCC;14'd7183:data <=32'h0004FFD3;14'd7184:data <=32'hFFFFFFDC;
14'd7185:data <=32'hFFFDFFE5;14'd7186:data <=32'hFFFFFFED;14'd7187:data <=32'h0005FFF2;
14'd7188:data <=32'h000DFFF4;14'd7189:data <=32'h0014FFF0;14'd7190:data <=32'h0018FFE9;
14'd7191:data <=32'h0019FFE0;14'd7192:data <=32'h0016FFD8;14'd7193:data <=32'h000FFFD1;
14'd7194:data <=32'h0005FFCD;14'd7195:data <=32'hFFFCFFCD;14'd7196:data <=32'hFFF3FFD0;
14'd7197:data <=32'hFFEBFFD4;14'd7198:data <=32'hFFE6FFDB;14'd7199:data <=32'hFFE3FFE1;
14'd7200:data <=32'hFFE1FFE8;14'd7201:data <=32'hFFE1FFEE;14'd7202:data <=32'hFFE3FFF4;
14'd7203:data <=32'hFFE6FFFA;14'd7204:data <=32'hFFEBFFFD;14'd7205:data <=32'hFFF2FFFF;
14'd7206:data <=32'hFFF8FFFE;14'd7207:data <=32'hFFFDFFF9;14'd7208:data <=32'h0000FFF3;
14'd7209:data <=32'h0000FFEB;14'd7210:data <=32'hFFFDFFE4;14'd7211:data <=32'hFFF6FFDF;
14'd7212:data <=32'hFFEDFFDC;14'd7213:data <=32'hFFE5FFDC;14'd7214:data <=32'hFFDDFFDF;
14'd7215:data <=32'hFFD7FFE3;14'd7216:data <=32'hFFD2FFE7;14'd7217:data <=32'hFFCEFFEB;
14'd7218:data <=32'hFFCBFFEF;14'd7219:data <=32'hFFC6FFF3;14'd7220:data <=32'hFFC0FFF8;
14'd7221:data <=32'hFFBAFFFF;14'd7222:data <=32'hFFB50008;14'd7223:data <=32'hFFB10013;
14'd7224:data <=32'hFFB00021;14'd7225:data <=32'hFFB1002E;14'd7226:data <=32'hFFB5003C;
14'd7227:data <=32'hFFBC004A;14'd7228:data <=32'hFFC50056;14'd7229:data <=32'hFFD00063;
14'd7230:data <=32'hFFDE006F;14'd7231:data <=32'hFFF00078;14'd7232:data <=32'h000C0020;
14'd7233:data <=32'h00080027;14'd7234:data <=32'h00050036;14'd7235:data <=32'h00140078;
14'd7236:data <=32'h003F0083;14'd7237:data <=32'h00570071;14'd7238:data <=32'h00690059;
14'd7239:data <=32'h0073003E;14'd7240:data <=32'h00750024;14'd7241:data <=32'h0072000D;
14'd7242:data <=32'h0069FFF8;14'd7243:data <=32'h005EFFE8;14'd7244:data <=32'h0050FFDB;
14'd7245:data <=32'h0042FFD2;14'd7246:data <=32'h0032FFCE;14'd7247:data <=32'h0023FFCD;
14'd7248:data <=32'h0015FFD2;14'd7249:data <=32'h000AFFD9;14'd7250:data <=32'h0004FFE3;
14'd7251:data <=32'h0003FFED;14'd7252:data <=32'h0006FFF5;14'd7253:data <=32'h000BFFFA;
14'd7254:data <=32'h0011FFFB;14'd7255:data <=32'h0016FFF9;14'd7256:data <=32'h0019FFF4;
14'd7257:data <=32'h0019FFEF;14'd7258:data <=32'h0018FFEB;14'd7259:data <=32'h0016FFE8;
14'd7260:data <=32'h0013FFE7;14'd7261:data <=32'h0011FFE6;14'd7262:data <=32'h0010FFE5;
14'd7263:data <=32'h000FFFE4;14'd7264:data <=32'h000DFFE2;14'd7265:data <=32'h000BFFE0;
14'd7266:data <=32'h0008FFDE;14'd7267:data <=32'h0005FFDE;14'd7268:data <=32'h0001FFDE;
14'd7269:data <=32'hFFFEFFDE;14'd7270:data <=32'hFFFCFFDE;14'd7271:data <=32'hFFFAFFDF;
14'd7272:data <=32'hFFF8FFDF;14'd7273:data <=32'hFFF5FFDF;14'd7274:data <=32'hFFF2FFDF;
14'd7275:data <=32'hFFEEFFE1;14'd7276:data <=32'hFFEBFFE3;14'd7277:data <=32'hFFE8FFE7;
14'd7278:data <=32'hFFE8FFEC;14'd7279:data <=32'hFFEAFFF0;14'd7280:data <=32'hFFEEFFF2;
14'd7281:data <=32'hFFF3FFF0;14'd7282:data <=32'hFFF7FFEC;14'd7283:data <=32'hFFF8FFE5;
14'd7284:data <=32'hFFF5FFDB;14'd7285:data <=32'hFFEDFFD3;14'd7286:data <=32'hFFE2FFCD;
14'd7287:data <=32'hFFD3FFCC;14'd7288:data <=32'hFFC4FFCE;14'd7289:data <=32'hFFB4FFD5;
14'd7290:data <=32'hFFA6FFE0;14'd7291:data <=32'hFF9AFFEE;14'd7292:data <=32'hFF910000;
14'd7293:data <=32'hFF8B0016;14'd7294:data <=32'hFF8A002F;14'd7295:data <=32'hFF900048;
14'd7296:data <=32'hFFC8002D;14'd7297:data <=32'hFFC5003D;14'd7298:data <=32'hFFC10048;
14'd7299:data <=32'hFFAC0058;14'd7300:data <=32'hFFD1007A;14'd7301:data <=32'hFFEA007C;
14'd7302:data <=32'h0001007A;14'd7303:data <=32'h00150071;14'd7304:data <=32'h00250066;
14'd7305:data <=32'h0031005A;14'd7306:data <=32'h003B004E;14'd7307:data <=32'h00420041;
14'd7308:data <=32'h00460034;14'd7309:data <=32'h00490027;14'd7310:data <=32'h0049001B;
14'd7311:data <=32'h0047000F;14'd7312:data <=32'h00420005;14'd7313:data <=32'h003CFFFD;
14'd7314:data <=32'h0036FFF8;14'd7315:data <=32'h0031FFF5;14'd7316:data <=32'h002DFFF2;
14'd7317:data <=32'h002AFFEF;14'd7318:data <=32'h0027FFEC;14'd7319:data <=32'h0023FFE8;
14'd7320:data <=32'h001DFFE5;14'd7321:data <=32'h0015FFE3;14'd7322:data <=32'h000DFFE4;
14'd7323:data <=32'h0006FFE8;14'd7324:data <=32'h0001FFEF;14'd7325:data <=32'h0000FFF7;
14'd7326:data <=32'h0002FFFE;14'd7327:data <=32'h00070005;14'd7328:data <=32'h000E0008;
14'd7329:data <=32'h00150007;14'd7330:data <=32'h001C0005;14'd7331:data <=32'h00220000;
14'd7332:data <=32'h0026FFF9;14'd7333:data <=32'h0028FFF2;14'd7334:data <=32'h0029FFE9;
14'd7335:data <=32'h0028FFE2;14'd7336:data <=32'h0024FFDA;14'd7337:data <=32'h001FFFD2;
14'd7338:data <=32'h0016FFCB;14'd7339:data <=32'h000CFFC8;14'd7340:data <=32'h0002FFC8;
14'd7341:data <=32'hFFF8FFCB;14'd7342:data <=32'hFFF0FFD1;14'd7343:data <=32'hFFECFFD9;
14'd7344:data <=32'hFFECFFE1;14'd7345:data <=32'hFFEFFFE7;14'd7346:data <=32'hFFF5FFE9;
14'd7347:data <=32'hFFFAFFE8;14'd7348:data <=32'hFFFEFFE3;14'd7349:data <=32'hFFFEFFDB;
14'd7350:data <=32'hFFFBFFD3;14'd7351:data <=32'hFFF4FFCC;14'd7352:data <=32'hFFEAFFC7;
14'd7353:data <=32'hFFDFFFC5;14'd7354:data <=32'hFFD3FFC5;14'd7355:data <=32'hFFC6FFC9;
14'd7356:data <=32'hFFBAFFCF;14'd7357:data <=32'hFFADFFD8;14'd7358:data <=32'hFFA2FFE4;
14'd7359:data <=32'hFF9AFFF5;14'd7360:data <=32'hFFA0FFD7;14'd7361:data <=32'hFF89FFEA;
14'd7362:data <=32'hFF82FFFE;14'd7363:data <=32'hFFA70007;14'd7364:data <=32'hFFBB0028;
14'd7365:data <=32'hFFC4002E;14'd7366:data <=32'hFFCD0031;14'd7367:data <=32'hFFD30032;
14'd7368:data <=32'hFFD70033;14'd7369:data <=32'hFFDA0035;14'd7370:data <=32'hFFDC0039;
14'd7371:data <=32'hFFE00040;14'd7372:data <=32'hFFE60046;14'd7373:data <=32'hFFEF004C;
14'd7374:data <=32'hFFFA0050;14'd7375:data <=32'h00050051;14'd7376:data <=32'h00120050;
14'd7377:data <=32'h001D004D;14'd7378:data <=32'h00290047;14'd7379:data <=32'h00330040;
14'd7380:data <=32'h003D0037;14'd7381:data <=32'h0046002A;14'd7382:data <=32'h004B001C;
14'd7383:data <=32'h004D000B;14'd7384:data <=32'h0049FFFB;14'd7385:data <=32'h0040FFEB;
14'd7386:data <=32'h0034FFE0;14'd7387:data <=32'h0024FFDA;14'd7388:data <=32'h0014FFDA;
14'd7389:data <=32'h0007FFDF;14'd7390:data <=32'hFFFDFFE8;14'd7391:data <=32'hFFF7FFF3;
14'd7392:data <=32'hFFF5FFFE;14'd7393:data <=32'hFFF80008;14'd7394:data <=32'hFFFD0010;
14'd7395:data <=32'h00040016;14'd7396:data <=32'h000C0019;14'd7397:data <=32'h0015001B;
14'd7398:data <=32'h001E001A;14'd7399:data <=32'h00270017;14'd7400:data <=32'h002F0010;
14'd7401:data <=32'h00360008;14'd7402:data <=32'h003AFFFD;14'd7403:data <=32'h003AFFF3;
14'd7404:data <=32'h0038FFE8;14'd7405:data <=32'h0034FFE0;14'd7406:data <=32'h002EFFD9;
14'd7407:data <=32'h0028FFD5;14'd7408:data <=32'h0023FFD2;14'd7409:data <=32'h0020FFD0;
14'd7410:data <=32'h001DFFCC;14'd7411:data <=32'h001AFFC7;14'd7412:data <=32'h0016FFC1;
14'd7413:data <=32'h0010FFBA;14'd7414:data <=32'h0005FFB4;14'd7415:data <=32'hFFFAFFB0;
14'd7416:data <=32'hFFEDFFB0;14'd7417:data <=32'hFFDFFFB3;14'd7418:data <=32'hFFD4FFB9;
14'd7419:data <=32'hFFCAFFC1;14'd7420:data <=32'hFFC2FFCA;14'd7421:data <=32'hFFBCFFD4;
14'd7422:data <=32'hFFB7FFDE;14'd7423:data <=32'hFFB5FFE9;14'd7424:data <=32'hFFE2FF9E;
14'd7425:data <=32'hFFC3FF9C;14'd7426:data <=32'hFFA9FFAC;14'd7427:data <=32'hFFBAFFF7;
14'd7428:data <=32'hFFD00014;14'd7429:data <=32'hFFDA0013;14'd7430:data <=32'hFFE2000F;
14'd7431:data <=32'hFFE60008;14'd7432:data <=32'hFFE50000;14'd7433:data <=32'hFFDFFFFB;
14'd7434:data <=32'hFFD6FFFA;14'd7435:data <=32'hFFCCFFFE;14'd7436:data <=32'hFFC40006;
14'd7437:data <=32'hFFBF0011;14'd7438:data <=32'hFFBE001E;14'd7439:data <=32'hFFC1002B;
14'd7440:data <=32'hFFC60038;14'd7441:data <=32'hFFCF0043;14'd7442:data <=32'hFFDA004D;
14'd7443:data <=32'hFFE80054;14'd7444:data <=32'hFFF80058;14'd7445:data <=32'h000A0059;
14'd7446:data <=32'h001B0054;14'd7447:data <=32'h002B004A;14'd7448:data <=32'h0037003C;
14'd7449:data <=32'h003E002B;14'd7450:data <=32'h003F001A;14'd7451:data <=32'h003B000A;
14'd7452:data <=32'h0033FFFE;14'd7453:data <=32'h0029FFF6;14'd7454:data <=32'h001FFFF3;
14'd7455:data <=32'h0016FFF2;14'd7456:data <=32'h000EFFF3;14'd7457:data <=32'h0008FFF6;
14'd7458:data <=32'h0003FFF9;14'd7459:data <=32'hFFFFFFFD;14'd7460:data <=32'hFFFC0003;
14'd7461:data <=32'hFFFA0008;14'd7462:data <=32'hFFFA000F;14'd7463:data <=32'hFFFC0017;
14'd7464:data <=32'h0000001E;14'd7465:data <=32'h00070024;14'd7466:data <=32'h000F0028;
14'd7467:data <=32'h00180029;14'd7468:data <=32'h00220029;14'd7469:data <=32'h002B0027;
14'd7470:data <=32'h00350023;14'd7471:data <=32'h003E001E;14'd7472:data <=32'h00480017;
14'd7473:data <=32'h0052000D;14'd7474:data <=32'h005B0000;14'd7475:data <=32'h0061FFEE;
14'd7476:data <=32'h0063FFDA;14'd7477:data <=32'h005FFFC4;14'd7478:data <=32'h0055FFAF;
14'd7479:data <=32'h0045FF9C;14'd7480:data <=32'h0030FF8F;14'd7481:data <=32'h0019FF87;
14'd7482:data <=32'h0001FF87;14'd7483:data <=32'hFFEAFF8C;14'd7484:data <=32'hFFD6FF95;
14'd7485:data <=32'hFFC6FFA2;14'd7486:data <=32'hFFB9FFB1;14'd7487:data <=32'hFFB1FFC3;
14'd7488:data <=32'h000BFFB8;14'd7489:data <=32'hFFFAFFAB;14'd7490:data <=32'hFFDFFFA5;
14'd7491:data <=32'hFFACFFCC;14'd7492:data <=32'hFFBEFFF2;14'd7493:data <=32'hFFC7FFFC;
14'd7494:data <=32'hFFD1FFFF;14'd7495:data <=32'hFFDAFFFF;14'd7496:data <=32'hFFDFFFFB;
14'd7497:data <=32'hFFE0FFF6;14'd7498:data <=32'hFFDCFFF3;14'd7499:data <=32'hFFD7FFF2;
14'd7500:data <=32'hFFD1FFF4;14'd7501:data <=32'hFFCCFFF9;14'd7502:data <=32'hFFC90000;
14'd7503:data <=32'hFFC70007;14'd7504:data <=32'hFFC7000F;14'd7505:data <=32'hFFC90016;
14'd7506:data <=32'hFFCB001E;14'd7507:data <=32'hFFCF0025;14'd7508:data <=32'hFFD5002D;
14'd7509:data <=32'hFFDC0032;14'd7510:data <=32'hFFE60037;14'd7511:data <=32'hFFF00038;
14'd7512:data <=32'hFFFA0037;14'd7513:data <=32'h00020033;14'd7514:data <=32'h0008002D;
14'd7515:data <=32'h000B0027;14'd7516:data <=32'h000C0022;14'd7517:data <=32'h000C001F;
14'd7518:data <=32'h000D001D;14'd7519:data <=32'h000E001C;14'd7520:data <=32'h0010001A;
14'd7521:data <=32'h00130017;14'd7522:data <=32'h00140013;14'd7523:data <=32'h0015000D;
14'd7524:data <=32'h00130007;14'd7525:data <=32'h000F0003;14'd7526:data <=32'h00080000;
14'd7527:data <=32'h00020000;14'd7528:data <=32'hFFFB0003;14'd7529:data <=32'hFFF50008;
14'd7530:data <=32'hFFF10010;14'd7531:data <=32'hFFF00018;14'd7532:data <=32'hFFF10022;
14'd7533:data <=32'hFFF5002C;14'd7534:data <=32'hFFFB0036;14'd7535:data <=32'h0005003F;
14'd7536:data <=32'h00130047;14'd7537:data <=32'h0024004B;14'd7538:data <=32'h0038004B;
14'd7539:data <=32'h004E0044;14'd7540:data <=32'h00610037;14'd7541:data <=32'h00710023;
14'd7542:data <=32'h007B000A;14'd7543:data <=32'h007DFFEF;14'd7544:data <=32'h0079FFD6;
14'd7545:data <=32'h006EFFBE;14'd7546:data <=32'h005EFFAC;14'd7547:data <=32'h004BFF9E;
14'd7548:data <=32'h0037FF95;14'd7549:data <=32'h0023FF90;14'd7550:data <=32'h000FFF90;
14'd7551:data <=32'hFFFCFF93;14'd7552:data <=32'h000FFFAF;14'd7553:data <=32'h0003FFA7;
14'd7554:data <=32'hFFF8FF9E;14'd7555:data <=32'hFFF3FF8E;14'd7556:data <=32'hFFF2FFAC;
14'd7557:data <=32'hFFEBFFB1;14'd7558:data <=32'hFFE4FFB5;14'd7559:data <=32'hFFDEFFB9;
14'd7560:data <=32'hFFD8FFBC;14'd7561:data <=32'hFFCFFFBF;14'd7562:data <=32'hFFC5FFC5;
14'd7563:data <=32'hFFBCFFCE;14'd7564:data <=32'hFFB4FFDA;14'd7565:data <=32'hFFB0FFE8;
14'd7566:data <=32'hFFB0FFF7;14'd7567:data <=32'hFFB40006;14'd7568:data <=32'hFFBB0011;
14'd7569:data <=32'hFFC5001A;14'd7570:data <=32'hFFCE001F;14'd7571:data <=32'hFFD80022;
14'd7572:data <=32'hFFE00022;14'd7573:data <=32'hFFE80021;14'd7574:data <=32'hFFEF001F;
14'd7575:data <=32'hFFF5001B;14'd7576:data <=32'hFFF90016;14'd7577:data <=32'hFFFB0010;
14'd7578:data <=32'hFFF90009;14'd7579:data <=32'hFFF50005;14'd7580:data <=32'hFFEF0003;
14'd7581:data <=32'hFFE90004;14'd7582:data <=32'hFFE4000A;14'd7583:data <=32'hFFE10011;
14'd7584:data <=32'hFFE30018;14'd7585:data <=32'hFFE7001F;14'd7586:data <=32'hFFEE0023;
14'd7587:data <=32'hFFF50024;14'd7588:data <=32'hFFFC0023;14'd7589:data <=32'h0001001F;
14'd7590:data <=32'h0003001A;14'd7591:data <=32'h00040016;14'd7592:data <=32'h00020012;
14'd7593:data <=32'hFFFF0010;14'd7594:data <=32'hFFFB0010;14'd7595:data <=32'hFFF80011;
14'd7596:data <=32'hFFF40013;14'd7597:data <=32'hFFF10018;14'd7598:data <=32'hFFEF001E;
14'd7599:data <=32'hFFEF0027;14'd7600:data <=32'hFFF10030;14'd7601:data <=32'hFFF7003A;
14'd7602:data <=32'h00010043;14'd7603:data <=32'h000F0049;14'd7604:data <=32'h001E004B;
14'd7605:data <=32'h002F0048;14'd7606:data <=32'h003E0040;14'd7607:data <=32'h004A0035;
14'd7608:data <=32'h00520027;14'd7609:data <=32'h00560019;14'd7610:data <=32'h0058000D;
14'd7611:data <=32'h00580002;14'd7612:data <=32'h0057FFF7;14'd7613:data <=32'h0056FFED;
14'd7614:data <=32'h0054FFE3;14'd7615:data <=32'h0051FFD8;14'd7616:data <=32'h0050FFB2;
14'd7617:data <=32'h0043FFA2;14'd7618:data <=32'h0039FF9E;14'd7619:data <=32'h0052FFC4;
14'd7620:data <=32'h0058FFD0;14'd7621:data <=32'h0054FFC1;14'd7622:data <=32'h004DFFB0;
14'd7623:data <=32'h0042FFA2;14'd7624:data <=32'h0033FF93;14'd7625:data <=32'h001EFF88;
14'd7626:data <=32'h0006FF82;14'd7627:data <=32'hFFECFF82;14'd7628:data <=32'hFFD2FF8A;
14'd7629:data <=32'hFFBCFF98;14'd7630:data <=32'hFFABFFAD;14'd7631:data <=32'hFFA2FFC4;
14'd7632:data <=32'hFF9EFFDB;14'd7633:data <=32'hFFA1FFF1;14'd7634:data <=32'hFFA90003;
14'd7635:data <=32'hFFB30012;14'd7636:data <=32'hFFC0001D;14'd7637:data <=32'hFFCE0024;
14'd7638:data <=32'hFFDC0027;14'd7639:data <=32'hFFEA0027;14'd7640:data <=32'hFFF70022;
14'd7641:data <=32'h0001001A;14'd7642:data <=32'h0007000F;14'd7643:data <=32'h00090003;
14'd7644:data <=32'h0006FFF9;14'd7645:data <=32'hFFFFFFF1;14'd7646:data <=32'hFFF6FFED;
14'd7647:data <=32'hFFEEFFED;14'd7648:data <=32'hFFE6FFF0;14'd7649:data <=32'hFFE1FFF5;
14'd7650:data <=32'hFFDFFFFA;14'd7651:data <=32'hFFDEFFFF;14'd7652:data <=32'hFFDD0003;
14'd7653:data <=32'hFFDD0006;14'd7654:data <=32'hFFDC0008;14'd7655:data <=32'hFFDA000C;
14'd7656:data <=32'hFFDA0010;14'd7657:data <=32'hFFD90015;14'd7658:data <=32'hFFDA001B;
14'd7659:data <=32'hFFDB0021;14'd7660:data <=32'hFFDF0026;14'd7661:data <=32'hFFE3002B;
14'd7662:data <=32'hFFE8002F;14'd7663:data <=32'hFFEC0032;14'd7664:data <=32'hFFF10035;
14'd7665:data <=32'hFFF80039;14'd7666:data <=32'hFFFE003A;14'd7667:data <=32'h0006003C;
14'd7668:data <=32'h000F003B;14'd7669:data <=32'h00180037;14'd7670:data <=32'h001E0031;
14'd7671:data <=32'h0022002A;14'd7672:data <=32'h00230023;14'd7673:data <=32'h0021001E;
14'd7674:data <=32'h001D001C;14'd7675:data <=32'h001B001E;14'd7676:data <=32'h001B0022;
14'd7677:data <=32'h001F0027;14'd7678:data <=32'h0026002B;14'd7679:data <=32'h0031002D;
14'd7680:data <=32'h0066000E;14'd7681:data <=32'h006DFFFD;14'd7682:data <=32'h0065FFF1;
14'd7683:data <=32'h0042001A;14'd7684:data <=32'h0057002A;14'd7685:data <=32'h0064001D;
14'd7686:data <=32'h006E000B;14'd7687:data <=32'h0075FFF7;14'd7688:data <=32'h0076FFDF;
14'd7689:data <=32'h0070FFC6;14'd7690:data <=32'h0064FFAE;14'd7691:data <=32'h0050FF9B;
14'd7692:data <=32'h0038FF8D;14'd7693:data <=32'h001EFF88;14'd7694:data <=32'h0005FF8A;
14'd7695:data <=32'hFFEFFF92;14'd7696:data <=32'hFFDDFF9E;14'd7697:data <=32'hFFD0FFAC;
14'd7698:data <=32'hFFC7FFBB;14'd7699:data <=32'hFFC2FFCA;14'd7700:data <=32'hFFBFFFD9;
14'd7701:data <=32'hFFC0FFE7;14'd7702:data <=32'hFFC3FFF4;14'd7703:data <=32'hFFC90000;
14'd7704:data <=32'hFFD20009;14'd7705:data <=32'hFFDC000E;14'd7706:data <=32'hFFE60010;
14'd7707:data <=32'hFFEF000F;14'd7708:data <=32'hFFF6000B;14'd7709:data <=32'hFFFB0007;
14'd7710:data <=32'hFFFD0002;14'd7711:data <=32'hFFFEFFFE;14'd7712:data <=32'hFFFFFFFB;
14'd7713:data <=32'h0000FFF7;14'd7714:data <=32'h0000FFF3;14'd7715:data <=32'h0000FFEE;
14'd7716:data <=32'hFFFEFFE7;14'd7717:data <=32'hFFF9FFE0;14'd7718:data <=32'hFFF1FFDB;
14'd7719:data <=32'hFFE6FFD7;14'd7720:data <=32'hFFDAFFD8;14'd7721:data <=32'hFFCDFFDC;
14'd7722:data <=32'hFFC2FFE4;14'd7723:data <=32'hFFB9FFF0;14'd7724:data <=32'hFFB3FFFE;
14'd7725:data <=32'hFFB2000D;14'd7726:data <=32'hFFB3001C;14'd7727:data <=32'hFFB8002A;
14'd7728:data <=32'hFFBF0036;14'd7729:data <=32'hFFCA0041;14'd7730:data <=32'hFFD7004A;
14'd7731:data <=32'hFFE5004F;14'd7732:data <=32'hFFF40050;14'd7733:data <=32'h0003004D;
14'd7734:data <=32'h00100045;14'd7735:data <=32'h0019003B;14'd7736:data <=32'h001D002F;
14'd7737:data <=32'h001C0024;14'd7738:data <=32'h0017001C;14'd7739:data <=32'h00100018;
14'd7740:data <=32'h0009001A;14'd7741:data <=32'h0005001F;14'd7742:data <=32'h00040027;
14'd7743:data <=32'h0007002F;14'd7744:data <=32'h0017003B;14'd7745:data <=32'h00220040;
14'd7746:data <=32'h002B0039;14'd7747:data <=32'h00200022;14'd7748:data <=32'h0030003A;
14'd7749:data <=32'h003B0036;14'd7750:data <=32'h0045002F;14'd7751:data <=32'h004E0026;
14'd7752:data <=32'h00560019;14'd7753:data <=32'h005B000A;14'd7754:data <=32'h005CFFF9;
14'd7755:data <=32'h0058FFE9;14'd7756:data <=32'h0050FFDB;14'd7757:data <=32'h0044FFD0;
14'd7758:data <=32'h0038FFCB;14'd7759:data <=32'h002DFFC8;14'd7760:data <=32'h0024FFC8;
14'd7761:data <=32'h001DFFC7;14'd7762:data <=32'h0017FFC8;14'd7763:data <=32'h0012FFC7;
14'd7764:data <=32'h000BFFC6;14'd7765:data <=32'h0004FFC6;14'd7766:data <=32'hFFFDFFC7;
14'd7767:data <=32'hFFF5FFCA;14'd7768:data <=32'hFFEEFFCE;14'd7769:data <=32'hFFE9FFD4;
14'd7770:data <=32'hFFE5FFDA;14'd7771:data <=32'hFFE3FFE0;14'd7772:data <=32'hFFE1FFE7;
14'd7773:data <=32'hFFE1FFED;14'd7774:data <=32'hFFE1FFF4;14'd7775:data <=32'hFFE3FFFB;
14'd7776:data <=32'hFFE80002;14'd7777:data <=32'hFFEF0008;14'd7778:data <=32'hFFF8000B;
14'd7779:data <=32'h00030009;14'd7780:data <=32'h000D0003;14'd7781:data <=32'h0015FFF9;
14'd7782:data <=32'h0017FFEC;14'd7783:data <=32'h0016FFDF;14'd7784:data <=32'h000FFFD1;
14'd7785:data <=32'h0003FFC8;14'd7786:data <=32'hFFF5FFC1;14'd7787:data <=32'hFFE5FFC0;
14'd7788:data <=32'hFFD6FFC3;14'd7789:data <=32'hFFC8FFC9;14'd7790:data <=32'hFFBDFFD3;
14'd7791:data <=32'hFFB2FFDE;14'd7792:data <=32'hFFACFFEC;14'd7793:data <=32'hFFA8FFFB;
14'd7794:data <=32'hFFA7000B;14'd7795:data <=32'hFFAB001B;14'd7796:data <=32'hFFB20029;
14'd7797:data <=32'hFFBC0034;14'd7798:data <=32'hFFC7003C;14'd7799:data <=32'hFFD4003F;
14'd7800:data <=32'hFFDF003F;14'd7801:data <=32'hFFE6003E;14'd7802:data <=32'hFFEB003C;
14'd7803:data <=32'hFFEE003B;14'd7804:data <=32'hFFF0003D;14'd7805:data <=32'hFFF30040;
14'd7806:data <=32'hFFF80044;14'd7807:data <=32'h00000048;14'd7808:data <=32'hFFF00013;
14'd7809:data <=32'hFFEA0020;14'd7810:data <=32'hFFF0002D;14'd7811:data <=32'h00200042;
14'd7812:data <=32'h00320053;14'd7813:data <=32'h003D0048;14'd7814:data <=32'h0045003B;
14'd7815:data <=32'h004A002E;14'd7816:data <=32'h004D001F;14'd7817:data <=32'h004D0011;
14'd7818:data <=32'h004A0003;14'd7819:data <=32'h0042FFF7;14'd7820:data <=32'h0038FFEF;
14'd7821:data <=32'h002DFFEB;14'd7822:data <=32'h0022FFEB;14'd7823:data <=32'h001AFFF0;
14'd7824:data <=32'h0017FFF7;14'd7825:data <=32'h0017FFFD;14'd7826:data <=32'h001C0001;
14'd7827:data <=32'h00220001;14'd7828:data <=32'h0027FFFE;14'd7829:data <=32'h002CFFF8;
14'd7830:data <=32'h002EFFF0;14'd7831:data <=32'h002DFFE8;14'd7832:data <=32'h002AFFE0;
14'd7833:data <=32'h0026FFDA;14'd7834:data <=32'h001FFFD4;14'd7835:data <=32'h0018FFCF;
14'd7836:data <=32'h000FFFCC;14'd7837:data <=32'h0006FFCC;14'd7838:data <=32'hFFFBFFCE;
14'd7839:data <=32'hFFF2FFD3;14'd7840:data <=32'hFFECFFDC;14'd7841:data <=32'hFFE8FFE6;
14'd7842:data <=32'hFFE9FFF1;14'd7843:data <=32'hFFEEFFFA;14'd7844:data <=32'hFFF60000;
14'd7845:data <=32'hFFFF0002;14'd7846:data <=32'h0008FFFF;14'd7847:data <=32'h000FFFF9;
14'd7848:data <=32'h0013FFF2;14'd7849:data <=32'h0014FFE9;14'd7850:data <=32'h0012FFE1;
14'd7851:data <=32'h000EFFDA;14'd7852:data <=32'h0009FFD5;14'd7853:data <=32'h0004FFD0;
14'd7854:data <=32'hFFFDFFCC;14'd7855:data <=32'hFFF6FFC9;14'd7856:data <=32'hFFEEFFC7;
14'd7857:data <=32'hFFE4FFC5;14'd7858:data <=32'hFFDAFFC7;14'd7859:data <=32'hFFD0FFCA;
14'd7860:data <=32'hFFC6FFCF;14'd7861:data <=32'hFFBEFFD6;14'd7862:data <=32'hFFB7FFDE;
14'd7863:data <=32'hFFB1FFE6;14'd7864:data <=32'hFFABFFEF;14'd7865:data <=32'hFFA6FFF9;
14'd7866:data <=32'hFFA00005;14'd7867:data <=32'hFF9C0013;14'd7868:data <=32'hFF9A0024;
14'd7869:data <=32'hFF9C0038;14'd7870:data <=32'hFFA3004D;14'd7871:data <=32'hFFB20060;
14'd7872:data <=32'hFFF20013;14'd7873:data <=32'hFFE80017;14'd7874:data <=32'hFFDC0024;
14'd7875:data <=32'hFFD50068;14'd7876:data <=32'hFFF30085;14'd7877:data <=32'h000D0080;
14'd7878:data <=32'h00230076;14'd7879:data <=32'h00350068;14'd7880:data <=32'h00440057;
14'd7881:data <=32'h004E0043;14'd7882:data <=32'h0053002E;14'd7883:data <=32'h0051001A;
14'd7884:data <=32'h004A0008;14'd7885:data <=32'h003FFFFA;14'd7886:data <=32'h0030FFF3;
14'd7887:data <=32'h0023FFF1;14'd7888:data <=32'h0017FFF5;14'd7889:data <=32'h0011FFFB;
14'd7890:data <=32'h000E0003;14'd7891:data <=32'h00100008;14'd7892:data <=32'h0014000C;
14'd7893:data <=32'h0018000E;14'd7894:data <=32'h001C000D;14'd7895:data <=32'h0020000B;
14'd7896:data <=32'h00230008;14'd7897:data <=32'h00250004;14'd7898:data <=32'h00280000;
14'd7899:data <=32'h0028FFFB;14'd7900:data <=32'h0029FFF5;14'd7901:data <=32'h0027FFEF;
14'd7902:data <=32'h0024FFE9;14'd7903:data <=32'h001FFFE5;14'd7904:data <=32'h0019FFE3;
14'd7905:data <=32'h0014FFE3;14'd7906:data <=32'h000FFFE5;14'd7907:data <=32'h000DFFE8;
14'd7908:data <=32'h000CFFEA;14'd7909:data <=32'h000DFFEB;14'd7910:data <=32'h000EFFEA;
14'd7911:data <=32'h000EFFE8;14'd7912:data <=32'h000CFFE6;14'd7913:data <=32'h000AFFE4;
14'd7914:data <=32'h0006FFE5;14'd7915:data <=32'h0004FFE6;14'd7916:data <=32'h0002FFE9;
14'd7917:data <=32'h0003FFEC;14'd7918:data <=32'h0006FFEE;14'd7919:data <=32'h000BFFEE;
14'd7920:data <=32'h000FFFEA;14'd7921:data <=32'h0013FFE5;14'd7922:data <=32'h0015FFDD;
14'd7923:data <=32'h0014FFD4;14'd7924:data <=32'h0011FFCA;14'd7925:data <=32'h000BFFC0;
14'd7926:data <=32'h0003FFB8;14'd7927:data <=32'hFFF7FFAF;14'd7928:data <=32'hFFE8FFA8;
14'd7929:data <=32'hFFD6FFA5;14'd7930:data <=32'hFFC1FFA6;14'd7931:data <=32'hFFAAFFAC;
14'd7932:data <=32'hFF94FFBA;14'd7933:data <=32'hFF81FFCF;14'd7934:data <=32'hFF74FFE9;
14'd7935:data <=32'hFF6F0008;14'd7936:data <=32'hFFBD0006;14'd7937:data <=32'hFFB4000F;
14'd7938:data <=32'hFFA90013;14'd7939:data <=32'hFF87001E;14'd7940:data <=32'hFF98004B;
14'd7941:data <=32'hFFAA0059;14'd7942:data <=32'hFFBD0063;14'd7943:data <=32'hFFD10068;
14'd7944:data <=32'hFFE4006A;14'd7945:data <=32'hFFF80067;14'd7946:data <=32'h00090061;
14'd7947:data <=32'h00170057;14'd7948:data <=32'h0021004A;14'd7949:data <=32'h0026003E;
14'd7950:data <=32'h00280033;14'd7951:data <=32'h0027002A;14'd7952:data <=32'h00260024;
14'd7953:data <=32'h00250020;14'd7954:data <=32'h0025001E;14'd7955:data <=32'h0027001A;
14'd7956:data <=32'h00290015;14'd7957:data <=32'h0029000F;14'd7958:data <=32'h00280008;
14'd7959:data <=32'h00250002;14'd7960:data <=32'h001FFFFE;14'd7961:data <=32'h001AFFFC;
14'd7962:data <=32'h0015FFFC;14'd7963:data <=32'h0011FFFE;14'd7964:data <=32'h000E0001;
14'd7965:data <=32'h000D0004;14'd7966:data <=32'h000D0006;14'd7967:data <=32'h000F0009;
14'd7968:data <=32'h0010000B;14'd7969:data <=32'h0013000E;14'd7970:data <=32'h0017000F;
14'd7971:data <=32'h001D0010;14'd7972:data <=32'h0023000E;14'd7973:data <=32'h002A0009;
14'd7974:data <=32'h002F0002;14'd7975:data <=32'h0032FFF9;14'd7976:data <=32'h0031FFEF;
14'd7977:data <=32'h002DFFE6;14'd7978:data <=32'h0025FFDF;14'd7979:data <=32'h001CFFDB;
14'd7980:data <=32'h0013FFDC;14'd7981:data <=32'h000DFFDF;14'd7982:data <=32'h0009FFE4;
14'd7983:data <=32'h0008FFEA;14'd7984:data <=32'h000BFFEE;14'd7985:data <=32'h000FFFF0;
14'd7986:data <=32'h0015FFF0;14'd7987:data <=32'h001AFFEC;14'd7988:data <=32'h001EFFE7;
14'd7989:data <=32'h0021FFE0;14'd7990:data <=32'h0023FFD6;14'd7991:data <=32'h0022FFCC;
14'd7992:data <=32'h001FFFBF;14'd7993:data <=32'h0017FFB2;14'd7994:data <=32'h000AFFA7;
14'd7995:data <=32'hFFF9FF9E;14'd7996:data <=32'hFFE4FF9A;14'd7997:data <=32'hFFCDFF9D;
14'd7998:data <=32'hFFB7FFA5;14'd7999:data <=32'hFFA5FFB4;14'd8000:data <=32'hFFBCFFAB;
14'd8001:data <=32'hFFA4FFB2;14'd8002:data <=32'hFF97FFBC;14'd8003:data <=32'hFFAFFFC8;
14'd8004:data <=32'hFFB0FFED;14'd8005:data <=32'hFFB0FFF6;14'd8006:data <=32'hFFB0FFFE;
14'd8007:data <=32'hFFB00006;14'd8008:data <=32'hFFB1000F;14'd8009:data <=32'hFFB30019;
14'd8010:data <=32'hFFB70022;14'd8011:data <=32'hFFBC002A;14'd8012:data <=32'hFFC10031;
14'd8013:data <=32'hFFC80038;14'd8014:data <=32'hFFCE003E;14'd8015:data <=32'hFFD50046;
14'd8016:data <=32'hFFDE004D;14'd8017:data <=32'hFFEA0053;14'd8018:data <=32'hFFF90057;
14'd8019:data <=32'h00090057;14'd8020:data <=32'h001A0052;14'd8021:data <=32'h002A0048;
14'd8022:data <=32'h00350039;14'd8023:data <=32'h003A0029;14'd8024:data <=32'h003B0018;
14'd8025:data <=32'h0037000A;14'd8026:data <=32'h002FFFFE;14'd8027:data <=32'h0025FFF6;
14'd8028:data <=32'h001BFFF2;14'd8029:data <=32'h0010FFF1;14'd8030:data <=32'h0006FFF3;
14'd8031:data <=32'hFFFEFFF7;14'd8032:data <=32'hFFF8FFFE;14'd8033:data <=32'hFFF40007;
14'd8034:data <=32'hFFF30011;14'd8035:data <=32'hFFF6001B;14'd8036:data <=32'hFFFC0024;
14'd8037:data <=32'h0006002A;14'd8038:data <=32'h0012002D;14'd8039:data <=32'h001D002B;
14'd8040:data <=32'h00270025;14'd8041:data <=32'h002E001D;14'd8042:data <=32'h00330015;
14'd8043:data <=32'h0034000C;14'd8044:data <=32'h00330006;14'd8045:data <=32'h00320001;
14'd8046:data <=32'h0032FFFD;14'd8047:data <=32'h0031FFFA;14'd8048:data <=32'h0033FFF7;
14'd8049:data <=32'h0034FFF2;14'd8050:data <=32'h0035FFEC;14'd8051:data <=32'h0036FFE6;
14'd8052:data <=32'h0034FFDE;14'd8053:data <=32'h0031FFD7;14'd8054:data <=32'h002EFFD0;
14'd8055:data <=32'h0029FFCA;14'd8056:data <=32'h0023FFC3;14'd8057:data <=32'h001DFFBD;
14'd8058:data <=32'h0015FFB7;14'd8059:data <=32'h000BFFB2;14'd8060:data <=32'hFFFEFFAF;
14'd8061:data <=32'hFFF1FFB0;14'd8062:data <=32'hFFE4FFB5;14'd8063:data <=32'hFFD9FFBD;
14'd8064:data <=32'h0018FF91;14'd8065:data <=32'hFFFEFF82;14'd8066:data <=32'hFFE4FF85;
14'd8067:data <=32'hFFDFFFCB;14'd8068:data <=32'hFFE4FFE7;14'd8069:data <=32'hFFE9FFE6;
14'd8070:data <=32'hFFEAFFE1;14'd8071:data <=32'hFFE9FFDC;14'd8072:data <=32'hFFE3FFD7;
14'd8073:data <=32'hFFDBFFD5;14'd8074:data <=32'hFFD3FFD5;14'd8075:data <=32'hFFC9FFD8;
14'd8076:data <=32'hFFBFFFDD;14'd8077:data <=32'hFFB5FFE5;14'd8078:data <=32'hFFACFFEF;
14'd8079:data <=32'hFFA5FFFE;14'd8080:data <=32'hFFA1000F;14'd8081:data <=32'hFFA30023;
14'd8082:data <=32'hFFAB0036;14'd8083:data <=32'hFFB80047;14'd8084:data <=32'hFFCA0054;
14'd8085:data <=32'hFFDF005A;14'd8086:data <=32'hFFF4005A;14'd8087:data <=32'h00060054;
14'd8088:data <=32'h0015004A;14'd8089:data <=32'h0020003D;14'd8090:data <=32'h0025002F;
14'd8091:data <=32'h00280023;14'd8092:data <=32'h00270017;14'd8093:data <=32'h0024000C;
14'd8094:data <=32'h001F0003;14'd8095:data <=32'h0018FFFC;14'd8096:data <=32'h000FFFF8;
14'd8097:data <=32'h0006FFF6;14'd8098:data <=32'hFFFCFFF7;14'd8099:data <=32'hFFF4FFFC;
14'd8100:data <=32'hFFEE0003;14'd8101:data <=32'hFFEB000C;14'd8102:data <=32'hFFEB0015;
14'd8103:data <=32'hFFED001C;14'd8104:data <=32'hFFF00023;14'd8105:data <=32'hFFF50028;
14'd8106:data <=32'hFFFA002D;14'd8107:data <=32'h00000032;14'd8108:data <=32'h00050036;
14'd8109:data <=32'h000E003B;14'd8110:data <=32'h0018003F;14'd8111:data <=32'h00250041;
14'd8112:data <=32'h00340040;14'd8113:data <=32'h0044003A;14'd8114:data <=32'h00520030;
14'd8115:data <=32'h005F0021;14'd8116:data <=32'h0067000F;14'd8117:data <=32'h006AFFFC;
14'd8118:data <=32'h0069FFE8;14'd8119:data <=32'h0063FFD5;14'd8120:data <=32'h005AFFC4;
14'd8121:data <=32'h004EFFB6;14'd8122:data <=32'h003FFFAA;14'd8123:data <=32'h002EFFA1;
14'd8124:data <=32'h001BFF9D;14'd8125:data <=32'h0007FF9E;14'd8126:data <=32'hFFF4FFA4;
14'd8127:data <=32'hFFE5FFAF;14'd8128:data <=32'h003BFFC9;14'd8129:data <=32'h0035FFB6;
14'd8130:data <=32'h0022FFA5;14'd8131:data <=32'hFFE6FFB9;14'd8132:data <=32'hFFE8FFDD;
14'd8133:data <=32'hFFEFFFE1;14'd8134:data <=32'hFFF3FFE1;14'd8135:data <=32'hFFF7FFDF;
14'd8136:data <=32'hFFF8FFDB;14'd8137:data <=32'hFFF6FFD7;14'd8138:data <=32'hFFF2FFD3;
14'd8139:data <=32'hFFEDFFD0;14'd8140:data <=32'hFFE6FFCE;14'd8141:data <=32'hFFDEFFCD;
14'd8142:data <=32'hFFD5FFCF;14'd8143:data <=32'hFFCAFFD2;14'd8144:data <=32'hFFC0FFDB;
14'd8145:data <=32'hFFB7FFE6;14'd8146:data <=32'hFFB2FFF4;14'd8147:data <=32'hFFB20003;
14'd8148:data <=32'hFFB60011;14'd8149:data <=32'hFFBE001D;14'd8150:data <=32'hFFC80025;
14'd8151:data <=32'hFFD3002A;14'd8152:data <=32'hFFDD002C;14'd8153:data <=32'hFFE4002B;
14'd8154:data <=32'hFFEB002A;14'd8155:data <=32'hFFF00029;14'd8156:data <=32'hFFF50028;
14'd8157:data <=32'hFFFA0026;14'd8158:data <=32'h00000024;14'd8159:data <=32'h00050020;
14'd8160:data <=32'h0008001B;14'd8161:data <=32'h000B0015;14'd8162:data <=32'h000B000F;
14'd8163:data <=32'h00090009;14'd8164:data <=32'h00050005;14'd8165:data <=32'h00010002;
14'd8166:data <=32'hFFFC0000;14'd8167:data <=32'hFFF7FFFF;14'd8168:data <=32'hFFF1FFFF;
14'd8169:data <=32'hFFEA0001;14'd8170:data <=32'hFFE30004;14'd8171:data <=32'hFFDB000B;
14'd8172:data <=32'hFFD50016;14'd8173:data <=32'hFFD10024;14'd8174:data <=32'hFFD30035;
14'd8175:data <=32'hFFD90046;14'd8176:data <=32'hFFE60056;14'd8177:data <=32'hFFF90062;
14'd8178:data <=32'h000F0069;14'd8179:data <=32'h00270069;14'd8180:data <=32'h003E0062;
14'd8181:data <=32'h00530056;14'd8182:data <=32'h00630046;14'd8183:data <=32'h00700032;
14'd8184:data <=32'h0077001C;14'd8185:data <=32'h007A0006;14'd8186:data <=32'h0078FFEF;
14'd8187:data <=32'h0072FFD9;14'd8188:data <=32'h0066FFC6;14'd8189:data <=32'h0056FFB7;
14'd8190:data <=32'h0042FFAD;14'd8191:data <=32'h002EFFA9;14'd8192:data <=32'h0033FFD1;
14'd8193:data <=32'h0030FFC9;14'd8194:data <=32'h002EFFBD;14'd8195:data <=32'h002EFFA7;
14'd8196:data <=32'h0026FFC1;14'd8197:data <=32'h0021FFBE;14'd8198:data <=32'h001BFFBA;
14'd8199:data <=32'h0015FFB6;14'd8200:data <=32'h000BFFB3;14'd8201:data <=32'h0000FFB2;
14'd8202:data <=32'hFFF4FFB4;14'd8203:data <=32'hFFEAFFB8;14'd8204:data <=32'hFFE1FFBE;
14'd8205:data <=32'hFFDAFFC5;14'd8206:data <=32'hFFD5FFCC;14'd8207:data <=32'hFFD0FFD4;
14'd8208:data <=32'hFFCCFFDD;14'd8209:data <=32'hFFCAFFE6;14'd8210:data <=32'hFFCAFFF0;
14'd8211:data <=32'hFFCCFFF9;14'd8212:data <=32'hFFD20002;14'd8213:data <=32'hFFDA0007;
14'd8214:data <=32'hFFE20008;14'd8215:data <=32'hFFE90007;14'd8216:data <=32'hFFED0002;
14'd8217:data <=32'hFFEEFFFD;14'd8218:data <=32'hFFEBFFF9;14'd8219:data <=32'hFFE7FFF8;
14'd8220:data <=32'hFFE2FFF9;14'd8221:data <=32'hFFDEFFFD;14'd8222:data <=32'hFFDC0002;
14'd8223:data <=32'hFFDC0008;14'd8224:data <=32'hFFDE000E;14'd8225:data <=32'hFFE10012;
14'd8226:data <=32'hFFE60015;14'd8227:data <=32'hFFEA0016;14'd8228:data <=32'hFFEF0016;
14'd8229:data <=32'hFFF30015;14'd8230:data <=32'hFFF60013;14'd8231:data <=32'hFFFA000F;
14'd8232:data <=32'hFFFB000A;14'd8233:data <=32'hFFF90004;14'd8234:data <=32'hFFF5FFFF;
14'd8235:data <=32'hFFEDFFFB;14'd8236:data <=32'hFFE4FFFB;14'd8237:data <=32'hFFD9FFFF;
14'd8238:data <=32'hFFD00008;14'd8239:data <=32'hFFC90015;14'd8240:data <=32'hFFC80024;
14'd8241:data <=32'hFFCB0034;14'd8242:data <=32'hFFD30043;14'd8243:data <=32'hFFDF004E;
14'd8244:data <=32'hFFEE0056;14'd8245:data <=32'hFFFD005A;14'd8246:data <=32'h000C005B;
14'd8247:data <=32'h001A0059;14'd8248:data <=32'h00290055;14'd8249:data <=32'h00360050;
14'd8250:data <=32'h00420047;14'd8251:data <=32'h004C003D;14'd8252:data <=32'h00550030;
14'd8253:data <=32'h005A0022;14'd8254:data <=32'h005C0015;14'd8255:data <=32'h005B0008;
14'd8256:data <=32'h005CFFE5;14'd8257:data <=32'h0057FFD9;14'd8258:data <=32'h0053FFD7;
14'd8259:data <=32'h00670000;14'd8260:data <=32'h006C000D;14'd8261:data <=32'h0073FFFA;
14'd8262:data <=32'h0075FFE4;14'd8263:data <=32'h0071FFCE;14'd8264:data <=32'h0067FFB8;
14'd8265:data <=32'h0056FFA5;14'd8266:data <=32'h0041FF97;14'd8267:data <=32'h002AFF8F;
14'd8268:data <=32'h0013FF8E;14'd8269:data <=32'hFFFEFF92;14'd8270:data <=32'hFFEAFF9A;
14'd8271:data <=32'hFFDAFFA5;14'd8272:data <=32'hFFCCFFB3;14'd8273:data <=32'hFFC3FFC3;
14'd8274:data <=32'hFFBEFFD6;14'd8275:data <=32'hFFBEFFE8;14'd8276:data <=32'hFFC4FFF9;
14'd8277:data <=32'hFFCE0006;14'd8278:data <=32'hFFDC000E;14'd8279:data <=32'hFFEA0011;
14'd8280:data <=32'hFFF6000E;14'd8281:data <=32'hFFFF0007;14'd8282:data <=32'h0004FFFE;
14'd8283:data <=32'h0005FFF5;14'd8284:data <=32'h0002FFEE;14'd8285:data <=32'hFFFDFFE9;
14'd8286:data <=32'hFFF7FFE6;14'd8287:data <=32'hFFF2FFE6;14'd8288:data <=32'hFFEDFFE6;
14'd8289:data <=32'hFFE9FFE8;14'd8290:data <=32'hFFE5FFEA;14'd8291:data <=32'hFFE2FFEC;
14'd8292:data <=32'hFFDFFFF0;14'd8293:data <=32'hFFDDFFF3;14'd8294:data <=32'hFFDBFFF7;
14'd8295:data <=32'hFFDBFFFB;14'd8296:data <=32'hFFDCFFFF;14'd8297:data <=32'hFFDD0001;
14'd8298:data <=32'hFFDD0002;14'd8299:data <=32'hFFDC0003;14'd8300:data <=32'hFFDA0004;
14'd8301:data <=32'hFFD70007;14'd8302:data <=32'hFFD4000A;14'd8303:data <=32'hFFD10011;
14'd8304:data <=32'hFFD10019;14'd8305:data <=32'hFFD40021;14'd8306:data <=32'hFFD90028;
14'd8307:data <=32'hFFE0002C;14'd8308:data <=32'hFFE7002E;14'd8309:data <=32'hFFEC002E;
14'd8310:data <=32'hFFF0002D;14'd8311:data <=32'hFFF1002C;14'd8312:data <=32'hFFF2002D;
14'd8313:data <=32'hFFF20030;14'd8314:data <=32'hFFF30034;14'd8315:data <=32'hFFF6003A;
14'd8316:data <=32'hFFFB003F;14'd8317:data <=32'h00000044;14'd8318:data <=32'h00080049;
14'd8319:data <=32'h0011004D;14'd8320:data <=32'h004C0039;14'd8321:data <=32'h00540031;
14'd8322:data <=32'h0050002A;14'd8323:data <=32'h0027004D;14'd8324:data <=32'h003A0067;
14'd8325:data <=32'h0052005F;14'd8326:data <=32'h0067004F;14'd8327:data <=32'h007A003A;
14'd8328:data <=32'h0085001F;14'd8329:data <=32'h00880003;14'd8330:data <=32'h0083FFE8;
14'd8331:data <=32'h0078FFD0;14'd8332:data <=32'h0069FFBC;14'd8333:data <=32'h0057FFAD;
14'd8334:data <=32'h0043FFA3;14'd8335:data <=32'h002EFF9D;14'd8336:data <=32'h0019FF9C;
14'd8337:data <=32'h0005FFA0;14'd8338:data <=32'hFFF3FFA8;14'd8339:data <=32'hFFE4FFB4;
14'd8340:data <=32'hFFDAFFC3;14'd8341:data <=32'hFFD6FFD3;14'd8342:data <=32'hFFD7FFE2;
14'd8343:data <=32'hFFDBFFEE;14'd8344:data <=32'hFFE2FFF7;14'd8345:data <=32'hFFEAFFFB;
14'd8346:data <=32'hFFF0FFFD;14'd8347:data <=32'hFFF5FFFD;14'd8348:data <=32'hFFF9FFFC;
14'd8349:data <=32'hFFFCFFFC;14'd8350:data <=32'hFFFFFFFB;14'd8351:data <=32'h0003FFFB;
14'd8352:data <=32'h0007FFF8;14'd8353:data <=32'h000AFFF4;14'd8354:data <=32'h000DFFEE;
14'd8355:data <=32'h000DFFE7;14'd8356:data <=32'h000BFFDF;14'd8357:data <=32'h0006FFD8;
14'd8358:data <=32'hFFFFFFD3;14'd8359:data <=32'hFFF7FFCF;14'd8360:data <=32'hFFEEFFCD;
14'd8361:data <=32'hFFE4FFCE;14'd8362:data <=32'hFFDBFFCF;14'd8363:data <=32'hFFD1FFD3;
14'd8364:data <=32'hFFC7FFD9;14'd8365:data <=32'hFFBFFFE1;14'd8366:data <=32'hFFB8FFED;
14'd8367:data <=32'hFFB3FFFB;14'd8368:data <=32'hFFB30009;14'd8369:data <=32'hFFB70018;
14'd8370:data <=32'hFFC00024;14'd8371:data <=32'hFFCB002D;14'd8372:data <=32'hFFD80031;
14'd8373:data <=32'hFFE4002F;14'd8374:data <=32'hFFED002B;14'd8375:data <=32'hFFF20024;
14'd8376:data <=32'hFFF3001E;14'd8377:data <=32'hFFF10018;14'd8378:data <=32'hFFED0016;
14'd8379:data <=32'hFFE80016;14'd8380:data <=32'hFFE30019;14'd8381:data <=32'hFFDE001F;
14'd8382:data <=32'hFFDB0027;14'd8383:data <=32'hFFDA0031;14'd8384:data <=32'hFFEE003F;
14'd8385:data <=32'hFFF2004B;14'd8386:data <=32'hFFF8004C;14'd8387:data <=32'hFFEF0039;
14'd8388:data <=32'hFFF7005C;14'd8389:data <=32'h00090062;14'd8390:data <=32'h001C0062;
14'd8391:data <=32'h002F005C;14'd8392:data <=32'h00400051;14'd8393:data <=32'h004C0043;
14'd8394:data <=32'h00540033;14'd8395:data <=32'h00570023;14'd8396:data <=32'h00570015;
14'd8397:data <=32'h00550008;14'd8398:data <=32'h0053FFFD;14'd8399:data <=32'h004FFFF2;
14'd8400:data <=32'h004AFFE8;14'd8401:data <=32'h0042FFDF;14'd8402:data <=32'h003BFFD8;
14'd8403:data <=32'h0031FFD3;14'd8404:data <=32'h0028FFD0;14'd8405:data <=32'h001FFFCF;
14'd8406:data <=32'h0018FFD0;14'd8407:data <=32'h0012FFD1;14'd8408:data <=32'h000DFFD2;
14'd8409:data <=32'h0008FFD3;14'd8410:data <=32'h0001FFD3;14'd8411:data <=32'hFFFAFFD6;
14'd8412:data <=32'hFFF3FFDA;14'd8413:data <=32'hFFEDFFE1;14'd8414:data <=32'hFFEAFFEB;
14'd8415:data <=32'hFFEAFFF5;14'd8416:data <=32'hFFEFFFFF;14'd8417:data <=32'hFFF70006;
14'd8418:data <=32'h0001000A;14'd8419:data <=32'h000C0009;14'd8420:data <=32'h00160004;
14'd8421:data <=32'h001EFFFC;14'd8422:data <=32'h0023FFF2;14'd8423:data <=32'h0025FFE6;
14'd8424:data <=32'h0023FFDB;14'd8425:data <=32'h001FFFCF;14'd8426:data <=32'h0017FFC4;
14'd8427:data <=32'h000CFFBB;14'd8428:data <=32'hFFFFFFB4;14'd8429:data <=32'hFFEFFFB1;
14'd8430:data <=32'hFFDEFFB3;14'd8431:data <=32'hFFCEFFB8;14'd8432:data <=32'hFFC0FFC3;
14'd8433:data <=32'hFFB6FFD1;14'd8434:data <=32'hFFB1FFE2;14'd8435:data <=32'hFFB1FFF1;
14'd8436:data <=32'hFFB5FFFE;14'd8437:data <=32'hFFBB0007;14'd8438:data <=32'hFFC1000D;
14'd8439:data <=32'hFFC70010;14'd8440:data <=32'hFFCA0012;14'd8441:data <=32'hFFCC0014;
14'd8442:data <=32'hFFCD0016;14'd8443:data <=32'hFFCD0019;14'd8444:data <=32'hFFCE001E;
14'd8445:data <=32'hFFCE0023;14'd8446:data <=32'hFFD00028;14'd8447:data <=32'hFFD2002D;
14'd8448:data <=32'hFFD9FFFC;14'd8449:data <=32'hFFC80005;14'd8450:data <=32'hFFC30015;
14'd8451:data <=32'hFFE60039;14'd8452:data <=32'hFFED0057;14'd8453:data <=32'hFFFC0058;
14'd8454:data <=32'h000B0055;14'd8455:data <=32'h0019004E;14'd8456:data <=32'h00240043;
14'd8457:data <=32'h002A0037;14'd8458:data <=32'h002B002B;14'd8459:data <=32'h00290021;
14'd8460:data <=32'h0024001B;14'd8461:data <=32'h00200017;14'd8462:data <=32'h001C0018;
14'd8463:data <=32'h001B0019;14'd8464:data <=32'h001D001B;14'd8465:data <=32'h0020001B;
14'd8466:data <=32'h0023001B;14'd8467:data <=32'h00280019;14'd8468:data <=32'h002C0017;
14'd8469:data <=32'h00310013;14'd8470:data <=32'h0036000E;14'd8471:data <=32'h003A0007;
14'd8472:data <=32'h003DFFFD;14'd8473:data <=32'h003EFFF2;14'd8474:data <=32'h003AFFE6;
14'd8475:data <=32'h0033FFDB;14'd8476:data <=32'h0027FFD3;14'd8477:data <=32'h001AFFCF;
14'd8478:data <=32'h000DFFD0;14'd8479:data <=32'h0001FFD5;14'd8480:data <=32'hFFF8FFDE;
14'd8481:data <=32'hFFF4FFE9;14'd8482:data <=32'hFFF4FFF3;14'd8483:data <=32'hFFF8FFFC;
14'd8484:data <=32'hFFFE0003;14'd8485:data <=32'h00060006;14'd8486:data <=32'h000E0007;
14'd8487:data <=32'h00150006;14'd8488:data <=32'h001C0002;14'd8489:data <=32'h0022FFFD;
14'd8490:data <=32'h0028FFF5;14'd8491:data <=32'h002BFFEC;14'd8492:data <=32'h002CFFE1;
14'd8493:data <=32'h0029FFD6;14'd8494:data <=32'h0024FFCB;14'd8495:data <=32'h001CFFC2;
14'd8496:data <=32'h0012FFBD;14'd8497:data <=32'h0007FFB9;14'd8498:data <=32'hFFFDFFB8;
14'd8499:data <=32'hFFF3FFB8;14'd8500:data <=32'hFFECFFB9;14'd8501:data <=32'hFFE4FFBA;
14'd8502:data <=32'hFFDBFFBA;14'd8503:data <=32'hFFD1FFBB;14'd8504:data <=32'hFFC5FFBD;
14'd8505:data <=32'hFFB7FFC2;14'd8506:data <=32'hFFAAFFCB;14'd8507:data <=32'hFF9EFFD9;
14'd8508:data <=32'hFF96FFE9;14'd8509:data <=32'hFF91FFFD;14'd8510:data <=32'hFF910010;
14'd8511:data <=32'hFF960023;14'd8512:data <=32'hFFEFFFF1;14'd8513:data <=32'hFFDEFFEB;
14'd8514:data <=32'hFFC7FFF2;14'd8515:data <=32'hFFA60036;14'd8516:data <=32'hFFB1005F;
14'd8517:data <=32'hFFC80069;14'd8518:data <=32'hFFE0006C;14'd8519:data <=32'hFFF80069;
14'd8520:data <=32'h000C005F;14'd8521:data <=32'h001C0050;14'd8522:data <=32'h0024003E;
14'd8523:data <=32'h0027002E;14'd8524:data <=32'h0023001F;14'd8525:data <=32'h001D0016;
14'd8526:data <=32'h00150011;14'd8527:data <=32'h000E0010;14'd8528:data <=32'h00080011;
14'd8529:data <=32'h00050014;14'd8530:data <=32'h00040018;14'd8531:data <=32'h0004001D;
14'd8532:data <=32'h00060021;14'd8533:data <=32'h000A0025;14'd8534:data <=32'h00100028;
14'd8535:data <=32'h0017002A;14'd8536:data <=32'h00200028;14'd8537:data <=32'h00290024;
14'd8538:data <=32'h0030001C;14'd8539:data <=32'h00340012;14'd8540:data <=32'h00340007;
14'd8541:data <=32'h0031FFFE;14'd8542:data <=32'h002BFFF7;14'd8543:data <=32'h0025FFF2;
14'd8544:data <=32'h001EFFF1;14'd8545:data <=32'h001AFFF2;14'd8546:data <=32'h0016FFF3;
14'd8547:data <=32'h0015FFF4;14'd8548:data <=32'h0014FFF5;14'd8549:data <=32'h0013FFF5;
14'd8550:data <=32'h0012FFF5;14'd8551:data <=32'h0010FFF6;14'd8552:data <=32'h000FFFF7;
14'd8553:data <=32'h000FFFF9;14'd8554:data <=32'h000FFFFC;14'd8555:data <=32'h0011FFFE;
14'd8556:data <=32'h00150000;14'd8557:data <=32'h0019FFFF;14'd8558:data <=32'h001EFFFE;
14'd8559:data <=32'h0023FFFC;14'd8560:data <=32'h0027FFF8;14'd8561:data <=32'h002CFFF3;
14'd8562:data <=32'h0030FFED;14'd8563:data <=32'h0035FFE5;14'd8564:data <=32'h0038FFDA;
14'd8565:data <=32'h003AFFCC;14'd8566:data <=32'h0037FFBC;14'd8567:data <=32'h0030FFAA;
14'd8568:data <=32'h0022FF99;14'd8569:data <=32'h000EFF8B;14'd8570:data <=32'hFFF6FF83;
14'd8571:data <=32'hFFDAFF81;14'd8572:data <=32'hFFBFFF88;14'd8573:data <=32'hFFA7FF95;
14'd8574:data <=32'hFF92FFA8;14'd8575:data <=32'hFF83FFBF;14'd8576:data <=32'hFFD5FFDE;
14'd8577:data <=32'hFFC9FFDA;14'd8578:data <=32'hFFB7FFD4;14'd8579:data <=32'hFF86FFD4;
14'd8580:data <=32'hFF7F0006;14'd8581:data <=32'hFF87001E;14'd8582:data <=32'hFF940032;
14'd8583:data <=32'hFFA60041;14'd8584:data <=32'hFFBA004A;14'd8585:data <=32'hFFCD004C;
14'd8586:data <=32'hFFDD004A;14'd8587:data <=32'hFFEA0044;14'd8588:data <=32'hFFF2003E;
14'd8589:data <=32'hFFF70038;14'd8590:data <=32'hFFFA0034;14'd8591:data <=32'hFFFD0032;
14'd8592:data <=32'h00010030;14'd8593:data <=32'h0005002D;14'd8594:data <=32'h0009002A;
14'd8595:data <=32'h000B0026;14'd8596:data <=32'h000D0022;14'd8597:data <=32'h000E001F;
14'd8598:data <=32'h000E001D;14'd8599:data <=32'h000E001C;14'd8600:data <=32'h000F001A;
14'd8601:data <=32'h00100019;14'd8602:data <=32'h00110016;14'd8603:data <=32'h00110013;
14'd8604:data <=32'h00100011;14'd8605:data <=32'h000E000F;14'd8606:data <=32'h000B000F;
14'd8607:data <=32'h00090011;14'd8608:data <=32'h00080015;14'd8609:data <=32'h000A0019;
14'd8610:data <=32'h000F001D;14'd8611:data <=32'h0016001E;14'd8612:data <=32'h001D001D;
14'd8613:data <=32'h00240018;14'd8614:data <=32'h00280012;14'd8615:data <=32'h002A000A;
14'd8616:data <=32'h00290003;14'd8617:data <=32'h0025FFFD;14'd8618:data <=32'h0021FFF9;
14'd8619:data <=32'h001CFFF8;14'd8620:data <=32'h0018FFF8;14'd8621:data <=32'h0015FFFA;
14'd8622:data <=32'h0013FFFD;14'd8623:data <=32'h00130000;14'd8624:data <=32'h00140005;
14'd8625:data <=32'h00170009;14'd8626:data <=32'h001E000C;14'd8627:data <=32'h0026000E;
14'd8628:data <=32'h0032000C;14'd8629:data <=32'h003E0006;14'd8630:data <=32'h0049FFFA;
14'd8631:data <=32'h0051FFEA;14'd8632:data <=32'h0054FFD6;14'd8633:data <=32'h0051FFC0;
14'd8634:data <=32'h0047FFAB;14'd8635:data <=32'h0036FF9A;14'd8636:data <=32'h0021FF8E;
14'd8637:data <=32'h000BFF88;14'd8638:data <=32'hFFF4FF87;14'd8639:data <=32'hFFDFFF8B;
14'd8640:data <=32'hFFF6FF98;14'd8641:data <=32'hFFE0FF8F;14'd8642:data <=32'hFFD1FF8C;
14'd8643:data <=32'hFFDBFF94;14'd8644:data <=32'hFFC6FFB6;14'd8645:data <=32'hFFBDFFC0;
14'd8646:data <=32'hFFB8FFCB;14'd8647:data <=32'hFFB4FFD7;14'd8648:data <=32'hFFB3FFE1;
14'd8649:data <=32'hFFB2FFE9;14'd8650:data <=32'hFFB2FFF1;14'd8651:data <=32'hFFB0FFF8;
14'd8652:data <=32'hFFAE0000;14'd8653:data <=32'hFFAC000A;14'd8654:data <=32'hFFAC0017;
14'd8655:data <=32'hFFAF0025;14'd8656:data <=32'hFFB70033;14'd8657:data <=32'hFFC2003F;
14'd8658:data <=32'hFFD10048;14'd8659:data <=32'hFFE1004C;14'd8660:data <=32'hFFF1004B;
14'd8661:data <=32'hFFFF0047;14'd8662:data <=32'h000A0040;14'd8663:data <=32'h00140037;
14'd8664:data <=32'h001B002D;14'd8665:data <=32'h001F0023;14'd8666:data <=32'h001F0017;
14'd8667:data <=32'h001E000C;14'd8668:data <=32'h00180002;14'd8669:data <=32'h0010FFFB;
14'd8670:data <=32'h0005FFF8;14'd8671:data <=32'hFFF9FFF8;14'd8672:data <=32'hFFEFFFFE;
14'd8673:data <=32'hFFE90007;14'd8674:data <=32'hFFE60013;14'd8675:data <=32'hFFE9001E;
14'd8676:data <=32'hFFEE0026;14'd8677:data <=32'hFFF7002D;14'd8678:data <=32'h0000002F;
14'd8679:data <=32'h0009002F;14'd8680:data <=32'h0010002D;14'd8681:data <=32'h00160029;
14'd8682:data <=32'h001A0026;14'd8683:data <=32'h001D0023;14'd8684:data <=32'h00200020;
14'd8685:data <=32'h0023001C;14'd8686:data <=32'h00250019;14'd8687:data <=32'h00270016;
14'd8688:data <=32'h00280014;14'd8689:data <=32'h00290012;14'd8690:data <=32'h002B0010;
14'd8691:data <=32'h002D000F;14'd8692:data <=32'h0032000E;14'd8693:data <=32'h0038000B;
14'd8694:data <=32'h003F0005;14'd8695:data <=32'h0045FFFD;14'd8696:data <=32'h0049FFF1;
14'd8697:data <=32'h0049FFE4;14'd8698:data <=32'h0045FFD7;14'd8699:data <=32'h003DFFCB;
14'd8700:data <=32'h0033FFC2;14'd8701:data <=32'h0029FFBD;14'd8702:data <=32'h001EFFBB;
14'd8703:data <=32'h0015FFBA;14'd8704:data <=32'h0055FFAA;14'd8705:data <=32'h0048FF8F;
14'd8706:data <=32'h0032FF82;14'd8707:data <=32'h0017FFBB;14'd8708:data <=32'h000DFFD2;
14'd8709:data <=32'h000CFFCF;14'd8710:data <=32'h000BFFCC;14'd8711:data <=32'h0009FFC7;
14'd8712:data <=32'h0005FFC1;14'd8713:data <=32'hFFFFFFBA;14'd8714:data <=32'hFFF6FFB3;
14'd8715:data <=32'hFFE9FFAE;14'd8716:data <=32'hFFD8FFAC;14'd8717:data <=32'hFFC6FFAF;
14'd8718:data <=32'hFFB3FFB9;14'd8719:data <=32'hFFA3FFC8;14'd8720:data <=32'hFF98FFDC;
14'd8721:data <=32'hFF94FFF4;14'd8722:data <=32'hFF96000A;14'd8723:data <=32'hFF9E001E;
14'd8724:data <=32'hFFAB002E;14'd8725:data <=32'hFFBA003A;14'd8726:data <=32'hFFCA0042;
14'd8727:data <=32'hFFDB0046;14'd8728:data <=32'hFFEB0046;14'd8729:data <=32'hFFFA0042;
14'd8730:data <=32'h0008003B;14'd8731:data <=32'h00130030;14'd8732:data <=32'h00190023;
14'd8733:data <=32'h001C0015;14'd8734:data <=32'h00190008;14'd8735:data <=32'h0012FFFD;
14'd8736:data <=32'h0008FFF6;14'd8737:data <=32'hFFFEFFF4;14'd8738:data <=32'hFFF4FFF5;
14'd8739:data <=32'hFFECFFF9;14'd8740:data <=32'hFFE7FFFF;14'd8741:data <=32'hFFE30005;
14'd8742:data <=32'hFFE1000A;14'd8743:data <=32'hFFE00010;14'd8744:data <=32'hFFDE0015;
14'd8745:data <=32'hFFDE001C;14'd8746:data <=32'hFFDE0024;14'd8747:data <=32'hFFE0002D;
14'd8748:data <=32'hFFE40037;14'd8749:data <=32'hFFEB003F;14'd8750:data <=32'hFFF50047;
14'd8751:data <=32'h0001004D;14'd8752:data <=32'h000E004F;14'd8753:data <=32'h001C004F;
14'd8754:data <=32'h002A004C;14'd8755:data <=32'h00370046;14'd8756:data <=32'h0043003F;
14'd8757:data <=32'h004F0035;14'd8758:data <=32'h00590027;14'd8759:data <=32'h00610017;
14'd8760:data <=32'h00640005;14'd8761:data <=32'h0062FFF2;14'd8762:data <=32'h005BFFE0;
14'd8763:data <=32'h004FFFD1;14'd8764:data <=32'h0040FFC7;14'd8765:data <=32'h0030FFC3;
14'd8766:data <=32'h0021FFC4;14'd8767:data <=32'h0015FFCA;14'd8768:data <=32'h005BFFFB;
14'd8769:data <=32'h0064FFE6;14'd8770:data <=32'h005DFFCC;14'd8771:data <=32'h001DFFC8;
14'd8772:data <=32'h0011FFE4;14'd8773:data <=32'h0014FFE7;14'd8774:data <=32'h0018FFE7;
14'd8775:data <=32'h001CFFE5;14'd8776:data <=32'h0021FFE0;14'd8777:data <=32'h0024FFD9;
14'd8778:data <=32'h0024FFCE;14'd8779:data <=32'h0020FFC2;14'd8780:data <=32'h0018FFB6;
14'd8781:data <=32'h000AFFAD;14'd8782:data <=32'hFFF9FFA8;14'd8783:data <=32'hFFE7FFA9;
14'd8784:data <=32'hFFD6FFAF;14'd8785:data <=32'hFFC8FFBA;14'd8786:data <=32'hFFBEFFC8;
14'd8787:data <=32'hFFB8FFD7;14'd8788:data <=32'hFFB6FFE5;14'd8789:data <=32'hFFB7FFF1;
14'd8790:data <=32'hFFBAFFFD;14'd8791:data <=32'hFFBE0007;14'd8792:data <=32'hFFC40010;
14'd8793:data <=32'hFFCA0018;14'd8794:data <=32'hFFD3001E;14'd8795:data <=32'hFFDD0022;
14'd8796:data <=32'hFFE60022;14'd8797:data <=32'hFFEF0021;14'd8798:data <=32'hFFF6001D;
14'd8799:data <=32'hFFFB0017;14'd8800:data <=32'hFFFE0012;14'd8801:data <=32'hFFFF000E;
14'd8802:data <=32'hFFFF000A;14'd8803:data <=32'hFFFF0006;14'd8804:data <=32'h00000002;
14'd8805:data <=32'hFFFFFFFD;14'd8806:data <=32'hFFFDFFF7;14'd8807:data <=32'hFFF8FFF1;
14'd8808:data <=32'hFFF0FFED;14'd8809:data <=32'hFFE5FFEB;14'd8810:data <=32'hFFD8FFEC;
14'd8811:data <=32'hFFCBFFF3;14'd8812:data <=32'hFFC0FFFE;14'd8813:data <=32'hFFB8000D;
14'd8814:data <=32'hFFB5001F;14'd8815:data <=32'hFFB70032;14'd8816:data <=32'hFFBE0044;
14'd8817:data <=32'hFFC90054;14'd8818:data <=32'hFFD80061;14'd8819:data <=32'hFFEB006C;
14'd8820:data <=32'hFFFF0072;14'd8821:data <=32'h00160073;14'd8822:data <=32'h002D0070;
14'd8823:data <=32'h00420066;14'd8824:data <=32'h00560056;14'd8825:data <=32'h00640042;
14'd8826:data <=32'h006C002B;14'd8827:data <=32'h006D0014;14'd8828:data <=32'h0067FFFE;
14'd8829:data <=32'h005DFFEE;14'd8830:data <=32'h0050FFE3;14'd8831:data <=32'h0043FFDD;
14'd8832:data <=32'h00390007;14'd8833:data <=32'h00400003;14'd8834:data <=32'h004AFFF5;
14'd8835:data <=32'h0051FFD8;14'd8836:data <=32'h0041FFEA;14'd8837:data <=32'h003EFFE5;
14'd8838:data <=32'h003AFFDF;14'd8839:data <=32'h0036FFDA;14'd8840:data <=32'h0032FFD5;
14'd8841:data <=32'h002EFFD1;14'd8842:data <=32'h002AFFCC;14'd8843:data <=32'h0025FFC6;
14'd8844:data <=32'h001DFFC0;14'd8845:data <=32'h0013FFBC;14'd8846:data <=32'h0008FFBA;
14'd8847:data <=32'hFFFCFFBC;14'd8848:data <=32'hFFF1FFC2;14'd8849:data <=32'hFFE9FFC9;
14'd8850:data <=32'hFFE4FFD3;14'd8851:data <=32'hFFE3FFDB;14'd8852:data <=32'hFFE5FFE2;
14'd8853:data <=32'hFFE8FFE6;14'd8854:data <=32'hFFEBFFE8;14'd8855:data <=32'hFFEBFFE8;
14'd8856:data <=32'hFFEBFFE8;14'd8857:data <=32'hFFE9FFE7;14'd8858:data <=32'hFFE7FFE9;
14'd8859:data <=32'hFFE5FFEB;14'd8860:data <=32'hFFE3FFED;14'd8861:data <=32'hFFE1FFF0;
14'd8862:data <=32'hFFE0FFF3;14'd8863:data <=32'hFFDFFFF6;14'd8864:data <=32'hFFDEFFFB;
14'd8865:data <=32'hFFDEFFFF;14'd8866:data <=32'hFFE00005;14'd8867:data <=32'hFFE4000A;
14'd8868:data <=32'hFFEA000D;14'd8869:data <=32'hFFF2000D;14'd8870:data <=32'hFFFA000B;
14'd8871:data <=32'hFFFF0004;14'd8872:data <=32'h0002FFFA;14'd8873:data <=32'hFFFFFFF0;
14'd8874:data <=32'hFFF9FFE7;14'd8875:data <=32'hFFEEFFE1;14'd8876:data <=32'hFFE1FFDF;
14'd8877:data <=32'hFFD4FFE1;14'd8878:data <=32'hFFC7FFE7;14'd8879:data <=32'hFFBDFFF2;
14'd8880:data <=32'hFFB5FFFF;14'd8881:data <=32'hFFB1000E;14'd8882:data <=32'hFFB0001D;
14'd8883:data <=32'hFFB2002D;14'd8884:data <=32'hFFB8003D;14'd8885:data <=32'hFFC1004C;
14'd8886:data <=32'hFFCF0058;14'd8887:data <=32'hFFDF0062;14'd8888:data <=32'hFFF10067;
14'd8889:data <=32'h00040067;14'd8890:data <=32'h00150062;14'd8891:data <=32'h0023005B;
14'd8892:data <=32'h002D0052;14'd8893:data <=32'h00340049;14'd8894:data <=32'h003A0041;
14'd8895:data <=32'h003E003B;14'd8896:data <=32'h00470017;14'd8897:data <=32'h00480012;
14'd8898:data <=32'h004B0012;14'd8899:data <=32'h0059003B;14'd8900:data <=32'h005B0046;
14'd8901:data <=32'h00670036;14'd8902:data <=32'h00700023;14'd8903:data <=32'h0074000E;
14'd8904:data <=32'h0073FFFA;14'd8905:data <=32'h006FFFE6;14'd8906:data <=32'h0067FFD4;
14'd8907:data <=32'h005CFFC3;14'd8908:data <=32'h004CFFB5;14'd8909:data <=32'h003AFFAB;
14'd8910:data <=32'h0026FFA5;14'd8911:data <=32'h0010FFA6;14'd8912:data <=32'hFFFDFFAD;
14'd8913:data <=32'hFFEDFFB9;14'd8914:data <=32'hFFE3FFC9;14'd8915:data <=32'hFFDFFFD9;
14'd8916:data <=32'hFFE1FFE7;14'd8917:data <=32'hFFE7FFF2;14'd8918:data <=32'hFFF0FFF9;
14'd8919:data <=32'hFFF8FFFB;14'd8920:data <=32'hFFFFFFFA;14'd8921:data <=32'h0005FFF8;
14'd8922:data <=32'h0008FFF4;14'd8923:data <=32'h000AFFEF;14'd8924:data <=32'h000BFFEA;
14'd8925:data <=32'h0009FFE5;14'd8926:data <=32'h0006FFE0;14'd8927:data <=32'h0002FFDC;
14'd8928:data <=32'hFFFBFFDA;14'd8929:data <=32'hFFF4FFDA;14'd8930:data <=32'hFFEEFFDC;
14'd8931:data <=32'hFFE9FFE1;14'd8932:data <=32'hFFE6FFE6;14'd8933:data <=32'hFFE6FFEC;
14'd8934:data <=32'hFFE8FFF0;14'd8935:data <=32'hFFEBFFF2;14'd8936:data <=32'hFFEEFFF1;
14'd8937:data <=32'hFFEFFFEE;14'd8938:data <=32'hFFEEFFEB;14'd8939:data <=32'hFFEAFFE8;
14'd8940:data <=32'hFFE5FFE7;14'd8941:data <=32'hFFDFFFE8;14'd8942:data <=32'hFFDAFFEA;
14'd8943:data <=32'hFFD6FFEF;14'd8944:data <=32'hFFD3FFF4;14'd8945:data <=32'hFFD1FFF8;
14'd8946:data <=32'hFFCFFFFC;14'd8947:data <=32'hFFCE0000;14'd8948:data <=32'hFFCC0004;
14'd8949:data <=32'hFFCB0009;14'd8950:data <=32'hFFC9000F;14'd8951:data <=32'hFFC90015;
14'd8952:data <=32'hFFCA001C;14'd8953:data <=32'hFFCB0022;14'd8954:data <=32'hFFCC0027;
14'd8955:data <=32'hFFCD002D;14'd8956:data <=32'hFFCE0034;14'd8957:data <=32'hFFCF003C;
14'd8958:data <=32'hFFD10048;14'd8959:data <=32'hFFD70055;14'd8960:data <=32'h001C0050;
14'd8961:data <=32'h0024004F;14'd8962:data <=32'h0024004D;14'd8963:data <=32'hFFF50067;
14'd8964:data <=32'h00000085;14'd8965:data <=32'h001B0085;14'd8966:data <=32'h0035007F;
14'd8967:data <=32'h004D0071;14'd8968:data <=32'h00600060;14'd8969:data <=32'h0070004B;
14'd8970:data <=32'h007A0034;14'd8971:data <=32'h007F001A;14'd8972:data <=32'h007E0000;
14'd8973:data <=32'h0077FFE8;14'd8974:data <=32'h006AFFD2;14'd8975:data <=32'h0057FFC1;
14'd8976:data <=32'h0042FFB7;14'd8977:data <=32'h002CFFB4;14'd8978:data <=32'h0018FFB7;
14'd8979:data <=32'h0009FFBF;14'd8980:data <=32'hFFFEFFCA;14'd8981:data <=32'hFFF8FFD5;
14'd8982:data <=32'hFFF6FFDF;14'd8983:data <=32'hFFF6FFE6;14'd8984:data <=32'hFFF7FFED;
14'd8985:data <=32'hFFF9FFF1;14'd8986:data <=32'hFFFBFFF6;14'd8987:data <=32'hFFFFFFFA;
14'd8988:data <=32'h0003FFFC;14'd8989:data <=32'h0007FFFD;14'd8990:data <=32'h000DFFFC;
14'd8991:data <=32'h0011FFFA;14'd8992:data <=32'h0014FFF6;14'd8993:data <=32'h0017FFF1;
14'd8994:data <=32'h0017FFEC;14'd8995:data <=32'h0016FFE8;14'd8996:data <=32'h0014FFE4;
14'd8997:data <=32'h0013FFE0;14'd8998:data <=32'h0012FFDB;14'd8999:data <=32'h000FFFD6;
14'd9000:data <=32'h000CFFD0;14'd9001:data <=32'h0005FFCA;14'd9002:data <=32'hFFFDFFC6;
14'd9003:data <=32'hFFF2FFC3;14'd9004:data <=32'hFFE6FFC4;14'd9005:data <=32'hFFDAFFC9;
14'd9006:data <=32'hFFD0FFD1;14'd9007:data <=32'hFFCAFFDC;14'd9008:data <=32'hFFC7FFE7;
14'd9009:data <=32'hFFC8FFF2;14'd9010:data <=32'hFFCCFFFA;14'd9011:data <=32'hFFD10000;
14'd9012:data <=32'hFFD70003;14'd9013:data <=32'hFFDC0004;14'd9014:data <=32'hFFDF0003;
14'd9015:data <=32'hFFE20001;14'd9016:data <=32'hFFE2FFFE;14'd9017:data <=32'hFFE1FFFA;
14'd9018:data <=32'hFFDDFFF7;14'd9019:data <=32'hFFD7FFF4;14'd9020:data <=32'hFFCDFFF4;
14'd9021:data <=32'hFFC1FFF8;14'd9022:data <=32'hFFB50000;14'd9023:data <=32'hFFAB000F;
14'd9024:data <=32'hFFC5002A;14'd9025:data <=32'hFFC20039;14'd9026:data <=32'hFFC5003F;
14'd9027:data <=32'hFFBE002C;14'd9028:data <=32'hFFBA0053;14'd9029:data <=32'hFFC90060;
14'd9030:data <=32'hFFDC0068;14'd9031:data <=32'hFFEF006C;14'd9032:data <=32'h0002006C;
14'd9033:data <=32'h00130069;14'd9034:data <=32'h00240063;14'd9035:data <=32'h0033005A;
14'd9036:data <=32'h0040004E;14'd9037:data <=32'h004A003F;14'd9038:data <=32'h0050002F;
14'd9039:data <=32'h0051001F;14'd9040:data <=32'h004F0011;14'd9041:data <=32'h00490005;
14'd9042:data <=32'h0043FFFC;14'd9043:data <=32'h003DFFF6;14'd9044:data <=32'h0037FFF2;
14'd9045:data <=32'h0033FFEE;14'd9046:data <=32'h0030FFEA;14'd9047:data <=32'h002CFFE5;
14'd9048:data <=32'h0026FFE0;14'd9049:data <=32'h001EFFDC;14'd9050:data <=32'h0015FFDB;
14'd9051:data <=32'h000BFFDC;14'd9052:data <=32'h0003FFE0;14'd9053:data <=32'hFFFDFFE7;
14'd9054:data <=32'hFFFAFFEF;14'd9055:data <=32'hFFFAFFF7;14'd9056:data <=32'hFFFCFFFF;
14'd9057:data <=32'h00000005;14'd9058:data <=32'h00060009;14'd9059:data <=32'h000D000C;
14'd9060:data <=32'h0016000D;14'd9061:data <=32'h001F000B;14'd9062:data <=32'h00280006;
14'd9063:data <=32'h0031FFFE;14'd9064:data <=32'h0037FFF3;14'd9065:data <=32'h003AFFE4;
14'd9066:data <=32'h0037FFD5;14'd9067:data <=32'h0030FFC6;14'd9068:data <=32'h0025FFBA;
14'd9069:data <=32'h0015FFB2;14'd9070:data <=32'h0005FFAF;14'd9071:data <=32'hFFF5FFB1;
14'd9072:data <=32'hFFE8FFB7;14'd9073:data <=32'hFFDEFFC0;14'd9074:data <=32'hFFD7FFC9;
14'd9075:data <=32'hFFD4FFD2;14'd9076:data <=32'hFFD3FFD9;14'd9077:data <=32'hFFD2FFE0;
14'd9078:data <=32'hFFD3FFE5;14'd9079:data <=32'hFFD4FFE9;14'd9080:data <=32'hFFD5FFEC;
14'd9081:data <=32'hFFD6FFEE;14'd9082:data <=32'hFFD6FFEE;14'd9083:data <=32'hFFD5FFED;
14'd9084:data <=32'hFFD2FFEC;14'd9085:data <=32'hFFCCFFEC;14'd9086:data <=32'hFFC3FFEE;
14'd9087:data <=32'hFFBAFFF4;14'd9088:data <=32'hFFD2FFD5;14'd9089:data <=32'hFFBAFFD9;
14'd9090:data <=32'hFFAEFFE8;14'd9091:data <=32'hFFC30013;14'd9092:data <=32'hFFBC0033;
14'd9093:data <=32'hFFC8003B;14'd9094:data <=32'hFFD5003F;14'd9095:data <=32'hFFE0003F;
14'd9096:data <=32'hFFE9003D;14'd9097:data <=32'hFFF0003A;14'd9098:data <=32'hFFF40037;
14'd9099:data <=32'hFFF90036;14'd9100:data <=32'hFFFC0034;14'd9101:data <=32'h00000033;
14'd9102:data <=32'h00030032;14'd9103:data <=32'h00050030;14'd9104:data <=32'h00070030;
14'd9105:data <=32'h00090031;14'd9106:data <=32'h000C0033;14'd9107:data <=32'h00120036;
14'd9108:data <=32'h001A0037;14'd9109:data <=32'h00240037;14'd9110:data <=32'h002F0032;
14'd9111:data <=32'h003A0029;14'd9112:data <=32'h0041001D;14'd9113:data <=32'h0044000D;
14'd9114:data <=32'h0042FFFF;14'd9115:data <=32'h003BFFF2;14'd9116:data <=32'h0032FFE9;
14'd9117:data <=32'h0026FFE3;14'd9118:data <=32'h001BFFE1;14'd9119:data <=32'h0010FFE3;
14'd9120:data <=32'h0007FFE7;14'd9121:data <=32'h0001FFED;14'd9122:data <=32'hFFFCFFF4;
14'd9123:data <=32'hFFFAFFFD;14'd9124:data <=32'hFFFA0006;14'd9125:data <=32'hFFFE0010;
14'd9126:data <=32'h00060017;14'd9127:data <=32'h0010001C;14'd9128:data <=32'h001D001C;
14'd9129:data <=32'h00280019;14'd9130:data <=32'h00330011;14'd9131:data <=32'h003B0006;
14'd9132:data <=32'h003EFFFA;14'd9133:data <=32'h003FFFED;14'd9134:data <=32'h003CFFE3;
14'd9135:data <=32'h0037FFDA;14'd9136:data <=32'h0031FFD2;14'd9137:data <=32'h002CFFCC;
14'd9138:data <=32'h0027FFC6;14'd9139:data <=32'h0022FFC0;14'd9140:data <=32'h001CFFBA;
14'd9141:data <=32'h0014FFB4;14'd9142:data <=32'h000AFFAE;14'd9143:data <=32'hFFFEFFAA;
14'd9144:data <=32'hFFF1FFA8;14'd9145:data <=32'hFFE4FFAA;14'd9146:data <=32'hFFD7FFAD;
14'd9147:data <=32'hFFCBFFB2;14'd9148:data <=32'hFFC0FFB9;14'd9149:data <=32'hFFB4FFC1;
14'd9150:data <=32'hFFA9FFCD;14'd9151:data <=32'hFFA0FFDA;14'd9152:data <=32'h0002FFD1;
14'd9153:data <=32'hFFEFFFC2;14'd9154:data <=32'hFFD5FFC1;14'd9155:data <=32'hFF9FFFFA;
14'd9156:data <=32'hFF990023;14'd9157:data <=32'hFFAA0033;14'd9158:data <=32'hFFBC003C;
14'd9159:data <=32'hFFCF003F;14'd9160:data <=32'hFFDF003C;14'd9161:data <=32'hFFEB0036;
14'd9162:data <=32'hFFF3002F;14'd9163:data <=32'hFFF80027;14'd9164:data <=32'hFFFA0020;
14'd9165:data <=32'hFFFA0019;14'd9166:data <=32'hFFF70015;14'd9167:data <=32'hFFF30011;
14'd9168:data <=32'hFFEE0011;14'd9169:data <=32'hFFE80013;14'd9170:data <=32'hFFE30019;
14'd9171:data <=32'hFFE10022;14'd9172:data <=32'hFFE3002C;14'd9173:data <=32'hFFE90036;
14'd9174:data <=32'hFFF4003E;14'd9175:data <=32'h00010041;14'd9176:data <=32'h000E0040;
14'd9177:data <=32'h001A003B;14'd9178:data <=32'h00230032;14'd9179:data <=32'h00290028;
14'd9180:data <=32'h002B001E;14'd9181:data <=32'h002B0015;14'd9182:data <=32'h0029000E;
14'd9183:data <=32'h00260008;14'd9184:data <=32'h00230003;14'd9185:data <=32'h001EFFFF;
14'd9186:data <=32'h001AFFFC;14'd9187:data <=32'h0014FFFB;14'd9188:data <=32'h000FFFFB;
14'd9189:data <=32'h000AFFFD;14'd9190:data <=32'h00070002;14'd9191:data <=32'h00060006;
14'd9192:data <=32'h0006000C;14'd9193:data <=32'h00090010;14'd9194:data <=32'h000C0013;
14'd9195:data <=32'h00110014;14'd9196:data <=32'h00150015;14'd9197:data <=32'h00180016;
14'd9198:data <=32'h001D0017;14'd9199:data <=32'h00220018;14'd9200:data <=32'h002A0019;
14'd9201:data <=32'h00330019;14'd9202:data <=32'h003E0015;14'd9203:data <=32'h004A000D;
14'd9204:data <=32'h00550000;14'd9205:data <=32'h005DFFEF;14'd9206:data <=32'h0060FFDB;
14'd9207:data <=32'h005EFFC5;14'd9208:data <=32'h0055FFB0;14'd9209:data <=32'h0048FF9D;
14'd9210:data <=32'h0036FF8E;14'd9211:data <=32'h0021FF82;14'd9212:data <=32'h0009FF7B;
14'd9213:data <=32'hFFF0FF79;14'd9214:data <=32'hFFD6FF7C;14'd9215:data <=32'hFFBCFF86;
14'd9216:data <=32'hFFFEFFCA;14'd9217:data <=32'hFFF4FFBD;14'd9218:data <=32'hFFE4FFAE;
14'd9219:data <=32'hFFADFF9E;14'd9220:data <=32'hFF93FFCA;14'd9221:data <=32'hFF94FFE2;
14'd9222:data <=32'hFF9AFFF6;14'd9223:data <=32'hFFA40006;14'd9224:data <=32'hFFAF0011;
14'd9225:data <=32'hFFBA0018;14'd9226:data <=32'hFFC4001C;14'd9227:data <=32'hFFCC001E;
14'd9228:data <=32'hFFD40020;14'd9229:data <=32'hFFDA001F;14'd9230:data <=32'hFFE0001F;
14'd9231:data <=32'hFFE4001D;14'd9232:data <=32'hFFE7001A;14'd9233:data <=32'hFFE80018;
14'd9234:data <=32'hFFE70017;14'd9235:data <=32'hFFE60019;14'd9236:data <=32'hFFE6001C;
14'd9237:data <=32'hFFE70020;14'd9238:data <=32'hFFEB0024;14'd9239:data <=32'hFFF10026;
14'd9240:data <=32'hFFF70026;14'd9241:data <=32'hFFFC0024;14'd9242:data <=32'h00000020;
14'd9243:data <=32'h0001001D;14'd9244:data <=32'h0000001A;14'd9245:data <=32'hFFFF0019;
14'd9246:data <=32'hFFFD001A;14'd9247:data <=32'hFFFE001C;14'd9248:data <=32'hFFFF001F;
14'd9249:data <=32'h00030021;14'd9250:data <=32'h00070022;14'd9251:data <=32'h000B0021;
14'd9252:data <=32'h000F001F;14'd9253:data <=32'h0012001C;14'd9254:data <=32'h00140019;
14'd9255:data <=32'h00150016;14'd9256:data <=32'h00150013;14'd9257:data <=32'h00150010;
14'd9258:data <=32'h0014000C;14'd9259:data <=32'h0012000A;14'd9260:data <=32'h000E0008;
14'd9261:data <=32'h00090009;14'd9262:data <=32'h0004000D;14'd9263:data <=32'h00010014;
14'd9264:data <=32'h0001001D;14'd9265:data <=32'h00050028;14'd9266:data <=32'h000F0031;
14'd9267:data <=32'h001D0038;14'd9268:data <=32'h002E003A;14'd9269:data <=32'h00410036;
14'd9270:data <=32'h0053002C;14'd9271:data <=32'h0061001C;14'd9272:data <=32'h006B0009;
14'd9273:data <=32'h0070FFF3;14'd9274:data <=32'h0070FFDD;14'd9275:data <=32'h006BFFC7;
14'd9276:data <=32'h0062FFB2;14'd9277:data <=32'h0054FF9F;14'd9278:data <=32'h0041FF8F;
14'd9279:data <=32'h002BFF84;14'd9280:data <=32'h0030FFA4;14'd9281:data <=32'h0021FF92;
14'd9282:data <=32'h0016FF86;14'd9283:data <=32'h001AFF89;14'd9284:data <=32'hFFF8FFA0;
14'd9285:data <=32'hFFEDFFA7;14'd9286:data <=32'hFFE5FFAD;14'd9287:data <=32'hFFDEFFB3;
14'd9288:data <=32'hFFD8FFB7;14'd9289:data <=32'hFFD0FFBB;14'd9290:data <=32'hFFC8FFC0;
14'd9291:data <=32'hFFBFFFC7;14'd9292:data <=32'hFFB7FFD1;14'd9293:data <=32'hFFB0FFDD;
14'd9294:data <=32'hFFADFFEA;14'd9295:data <=32'hFFADFFF8;14'd9296:data <=32'hFFB00005;
14'd9297:data <=32'hFFB40010;14'd9298:data <=32'hFFBB001A;14'd9299:data <=32'hFFC20024;
14'd9300:data <=32'hFFCB002B;14'd9301:data <=32'hFFD60031;14'd9302:data <=32'hFFE30035;
14'd9303:data <=32'hFFF00034;14'd9304:data <=32'hFFFD002F;14'd9305:data <=32'h00070026;
14'd9306:data <=32'h000D001B;14'd9307:data <=32'h000E000F;14'd9308:data <=32'h000A0005;
14'd9309:data <=32'h0003FFFD;14'd9310:data <=32'hFFF9FFF9;14'd9311:data <=32'hFFF0FFFA;
14'd9312:data <=32'hFFE8FFFF;14'd9313:data <=32'hFFE30005;14'd9314:data <=32'hFFE1000C;
14'd9315:data <=32'hFFE00014;14'd9316:data <=32'hFFE3001A;14'd9317:data <=32'hFFE60020;
14'd9318:data <=32'hFFEA0025;14'd9319:data <=32'hFFEF0029;14'd9320:data <=32'hFFF5002B;
14'd9321:data <=32'hFFFC002C;14'd9322:data <=32'h0002002B;14'd9323:data <=32'h00070028;
14'd9324:data <=32'h000A0025;14'd9325:data <=32'h000B0020;14'd9326:data <=32'h000A001E;
14'd9327:data <=32'h0008001E;14'd9328:data <=32'h00060020;14'd9329:data <=32'h00050025;
14'd9330:data <=32'h0007002B;14'd9331:data <=32'h000E0032;14'd9332:data <=32'h00170036;
14'd9333:data <=32'h00220037;14'd9334:data <=32'h002F0035;14'd9335:data <=32'h003A002F;
14'd9336:data <=32'h00430026;14'd9337:data <=32'h0049001C;14'd9338:data <=32'h004E0011;
14'd9339:data <=32'h00500007;14'd9340:data <=32'h0051FFFB;14'd9341:data <=32'h0051FFF0;
14'd9342:data <=32'h004FFFE5;14'd9343:data <=32'h004BFFDA;14'd9344:data <=32'h007CFFDD;
14'd9345:data <=32'h007BFFBE;14'd9346:data <=32'h006DFFAB;14'd9347:data <=32'h0046FFD5;
14'd9348:data <=32'h0033FFE5;14'd9349:data <=32'h0035FFE1;14'd9350:data <=32'h0038FFDB;
14'd9351:data <=32'h003BFFD1;14'd9352:data <=32'h003AFFC4;14'd9353:data <=32'h0035FFB5;
14'd9354:data <=32'h002AFFA6;14'd9355:data <=32'h001AFF9B;14'd9356:data <=32'h0006FF94;
14'd9357:data <=32'hFFF1FF92;14'd9358:data <=32'hFFDBFF97;14'd9359:data <=32'hFFC8FFA1;
14'd9360:data <=32'hFFB8FFAE;14'd9361:data <=32'hFFACFFBF;14'd9362:data <=32'hFFA4FFD1;
14'd9363:data <=32'hFF9FFFE4;14'd9364:data <=32'hFF9FFFF8;14'd9365:data <=32'hFFA5000C;
14'd9366:data <=32'hFFAF001D;14'd9367:data <=32'hFFBE002B;14'd9368:data <=32'hFFD00033;
14'd9369:data <=32'hFFE20035;14'd9370:data <=32'hFFF40031;14'd9371:data <=32'h00010029;
14'd9372:data <=32'h0009001D;14'd9373:data <=32'h000D0010;14'd9374:data <=32'h000C0005;
14'd9375:data <=32'h0008FFFC;14'd9376:data <=32'h0002FFF6;14'd9377:data <=32'hFFFCFFF2;
14'd9378:data <=32'hFFF5FFF0;14'd9379:data <=32'hFFEFFFF0;14'd9380:data <=32'hFFE9FFF0;
14'd9381:data <=32'hFFE3FFF2;14'd9382:data <=32'hFFDCFFF5;14'd9383:data <=32'hFFD6FFFA;
14'd9384:data <=32'hFFD10001;14'd9385:data <=32'hFFCE0009;14'd9386:data <=32'hFFCD0012;
14'd9387:data <=32'hFFCD001B;14'd9388:data <=32'hFFD00023;14'd9389:data <=32'hFFD3002B;
14'd9390:data <=32'hFFD70032;14'd9391:data <=32'hFFDC0039;14'd9392:data <=32'hFFE20040;
14'd9393:data <=32'hFFE90048;14'd9394:data <=32'hFFF4004F;14'd9395:data <=32'h00010054;
14'd9396:data <=32'h00100056;14'd9397:data <=32'h00200054;14'd9398:data <=32'h002F004C;
14'd9399:data <=32'h003C0041;14'd9400:data <=32'h00450033;14'd9401:data <=32'h00480024;
14'd9402:data <=32'h00470016;14'd9403:data <=32'h0044000B;14'd9404:data <=32'h003F0003;
14'd9405:data <=32'h0038FFFD;14'd9406:data <=32'h0033FFF9;14'd9407:data <=32'h002EFFF7;
14'd9408:data <=32'h005C0034;14'd9409:data <=32'h006E0023;14'd9410:data <=32'h00710009;
14'd9411:data <=32'h0032FFF3;14'd9412:data <=32'h001F000A;14'd9413:data <=32'h0025000E;
14'd9414:data <=32'h002F0010;14'd9415:data <=32'h003A000D;14'd9416:data <=32'h00460005;
14'd9417:data <=32'h004FFFF7;14'd9418:data <=32'h0053FFE6;14'd9419:data <=32'h0051FFD3;
14'd9420:data <=32'h004AFFC1;14'd9421:data <=32'h003DFFB3;14'd9422:data <=32'h002DFFA9;
14'd9423:data <=32'h001CFFA2;14'd9424:data <=32'h000BFFA0;14'd9425:data <=32'hFFFAFFA1;
14'd9426:data <=32'hFFEAFFA5;14'd9427:data <=32'hFFDBFFAD;14'd9428:data <=32'hFFCEFFB8;
14'd9429:data <=32'hFFC4FFC5;14'd9430:data <=32'hFFBEFFD5;14'd9431:data <=32'hFFBCFFE5;
14'd9432:data <=32'hFFBFFFF4;14'd9433:data <=32'hFFC60000;14'd9434:data <=32'hFFCF0009;
14'd9435:data <=32'hFFD9000D;14'd9436:data <=32'hFFE1000F;14'd9437:data <=32'hFFE8000F;
14'd9438:data <=32'hFFED000E;14'd9439:data <=32'hFFF2000C;14'd9440:data <=32'hFFF6000C;
14'd9441:data <=32'hFFFA0009;14'd9442:data <=32'hFFFF0007;14'd9443:data <=32'h00030002;
14'd9444:data <=32'h0007FFFB;14'd9445:data <=32'h0007FFF2;14'd9446:data <=32'h0004FFE9;
14'd9447:data <=32'hFFFEFFE1;14'd9448:data <=32'hFFF5FFDA;14'd9449:data <=32'hFFEAFFD7;
14'd9450:data <=32'hFFDDFFD6;14'd9451:data <=32'hFFD0FFD9;14'd9452:data <=32'hFFC4FFDF;
14'd9453:data <=32'hFFB8FFE8;14'd9454:data <=32'hFFAFFFF4;14'd9455:data <=32'hFFA70003;
14'd9456:data <=32'hFFA30015;14'd9457:data <=32'hFFA30029;14'd9458:data <=32'hFFA8003E;
14'd9459:data <=32'hFFB30051;14'd9460:data <=32'hFFC40062;14'd9461:data <=32'hFFD9006E;
14'd9462:data <=32'hFFF10073;14'd9463:data <=32'h00090071;14'd9464:data <=32'h001E0069;
14'd9465:data <=32'h002F005C;14'd9466:data <=32'h003A004C;14'd9467:data <=32'h0040003D;
14'd9468:data <=32'h0042002E;14'd9469:data <=32'h00410021;14'd9470:data <=32'h003E0017;
14'd9471:data <=32'h003A000E;14'd9472:data <=32'h00230031;14'd9473:data <=32'h002D0031;
14'd9474:data <=32'h003B0029;14'd9475:data <=32'h0047000A;14'd9476:data <=32'h00310019;
14'd9477:data <=32'h00320018;14'd9478:data <=32'h00360017;14'd9479:data <=32'h003A0014;
14'd9480:data <=32'h0041000F;14'd9481:data <=32'h00470006;14'd9482:data <=32'h004AFFFB;
14'd9483:data <=32'h0049FFEE;14'd9484:data <=32'h0044FFE2;14'd9485:data <=32'h003CFFD8;
14'd9486:data <=32'h0033FFD2;14'd9487:data <=32'h0029FFCE;14'd9488:data <=32'h0021FFCD;
14'd9489:data <=32'h001AFFCD;14'd9490:data <=32'h0014FFCD;14'd9491:data <=32'h000EFFCE;
14'd9492:data <=32'h0009FFCF;14'd9493:data <=32'h0003FFD1;14'd9494:data <=32'hFFFFFFD3;
14'd9495:data <=32'hFFFBFFD6;14'd9496:data <=32'hFFF8FFD9;14'd9497:data <=32'hFFF7FFDC;
14'd9498:data <=32'hFFF6FFDD;14'd9499:data <=32'hFFF5FFDE;14'd9500:data <=32'hFFF2FFDE;
14'd9501:data <=32'hFFEEFFDF;14'd9502:data <=32'hFFE9FFE1;14'd9503:data <=32'hFFE4FFE5;
14'd9504:data <=32'hFFE1FFEC;14'd9505:data <=32'hFFE0FFF5;14'd9506:data <=32'hFFE3FFFD;
14'd9507:data <=32'hFFEA0004;14'd9508:data <=32'hFFF30007;14'd9509:data <=32'hFFFC0006;
14'd9510:data <=32'h00050002;14'd9511:data <=32'h000BFFFA;14'd9512:data <=32'h000DFFF0;
14'd9513:data <=32'h000DFFE6;14'd9514:data <=32'h0009FFDC;14'd9515:data <=32'h0002FFD3;
14'd9516:data <=32'hFFF7FFCC;14'd9517:data <=32'hFFEBFFC7;14'd9518:data <=32'hFFDDFFC5;
14'd9519:data <=32'hFFCDFFC6;14'd9520:data <=32'hFFBDFFCC;14'd9521:data <=32'hFFAEFFD7;
14'd9522:data <=32'hFFA2FFE7;14'd9523:data <=32'hFF9BFFFB;14'd9524:data <=32'hFF99000F;
14'd9525:data <=32'hFF9D0024;14'd9526:data <=32'hFFA60036;14'd9527:data <=32'hFFB30044;
14'd9528:data <=32'hFFC1004D;14'd9529:data <=32'hFFD00053;14'd9530:data <=32'hFFDC0055;
14'd9531:data <=32'hFFE80055;14'd9532:data <=32'hFFF20056;14'd9533:data <=32'hFFFC0056;
14'd9534:data <=32'h00060055;14'd9535:data <=32'h00100053;14'd9536:data <=32'h00230030;
14'd9537:data <=32'h0024002D;14'd9538:data <=32'h00260030;14'd9539:data <=32'h00290059;
14'd9540:data <=32'h00220065;14'd9541:data <=32'h00320060;14'd9542:data <=32'h00410058;
14'd9543:data <=32'h004F004C;14'd9544:data <=32'h005C003E;14'd9545:data <=32'h0065002B;
14'd9546:data <=32'h006A0016;14'd9547:data <=32'h00680000;14'd9548:data <=32'h0060FFEB;
14'd9549:data <=32'h0052FFDB;14'd9550:data <=32'h0042FFD0;14'd9551:data <=32'h0031FFCC;
14'd9552:data <=32'h0021FFCC;14'd9553:data <=32'h0015FFD1;14'd9554:data <=32'h000CFFD8;
14'd9555:data <=32'h0006FFDF;14'd9556:data <=32'h0003FFE7;14'd9557:data <=32'h0003FFEE;
14'd9558:data <=32'h0004FFF3;14'd9559:data <=32'h0007FFF8;14'd9560:data <=32'h000CFFFB;
14'd9561:data <=32'h0012FFFB;14'd9562:data <=32'h0018FFF9;14'd9563:data <=32'h001DFFF4;
14'd9564:data <=32'h001FFFEC;14'd9565:data <=32'h001EFFE3;14'd9566:data <=32'h0019FFDC;
14'd9567:data <=32'h0011FFD7;14'd9568:data <=32'h0008FFD5;14'd9569:data <=32'h0000FFD7;
14'd9570:data <=32'hFFFAFFDB;14'd9571:data <=32'hFFF6FFE1;14'd9572:data <=32'hFFF6FFE7;
14'd9573:data <=32'hFFF7FFEB;14'd9574:data <=32'hFFFAFFEE;14'd9575:data <=32'hFFFEFFEE;
14'd9576:data <=32'h0000FFED;14'd9577:data <=32'h0002FFEA;14'd9578:data <=32'h0002FFE7;
14'd9579:data <=32'h0002FFE3;14'd9580:data <=32'h0000FFE0;14'd9581:data <=32'hFFFEFFDC;
14'd9582:data <=32'hFFFBFFD8;14'd9583:data <=32'hFFF6FFD4;14'd9584:data <=32'hFFEFFFD1;
14'd9585:data <=32'hFFE7FFD0;14'd9586:data <=32'hFFDFFFD1;14'd9587:data <=32'hFFD6FFD4;
14'd9588:data <=32'hFFCEFFD9;14'd9589:data <=32'hFFC9FFE0;14'd9590:data <=32'hFFC5FFE6;
14'd9591:data <=32'hFFC2FFEC;14'd9592:data <=32'hFFC0FFF0;14'd9593:data <=32'hFFBCFFF4;
14'd9594:data <=32'hFFB7FFF9;14'd9595:data <=32'hFFB00000;14'd9596:data <=32'hFFAA000B;
14'd9597:data <=32'hFFA40018;14'd9598:data <=32'hFFA20029;14'd9599:data <=32'hFFA5003C;
14'd9600:data <=32'hFFF20049;14'd9601:data <=32'hFFF80049;14'd9602:data <=32'hFFF50046;
14'd9603:data <=32'hFFBC0053;14'd9604:data <=32'hFFB70073;14'd9605:data <=32'hFFCE0081;
14'd9606:data <=32'hFFE7008A;14'd9607:data <=32'h0002008D;14'd9608:data <=32'h001F0089;
14'd9609:data <=32'h003A007E;14'd9610:data <=32'h0051006C;14'd9611:data <=32'h00620054;
14'd9612:data <=32'h006B003A;14'd9613:data <=32'h006C0020;14'd9614:data <=32'h00650008;
14'd9615:data <=32'h005AFFF5;14'd9616:data <=32'h004CFFE8;14'd9617:data <=32'h003EFFE1;
14'd9618:data <=32'h0030FFDD;14'd9619:data <=32'h0024FFDD;14'd9620:data <=32'h0019FFDF;
14'd9621:data <=32'h0010FFE3;14'd9622:data <=32'h000AFFE8;14'd9623:data <=32'h0005FFEE;
14'd9624:data <=32'h0003FFF6;14'd9625:data <=32'h0003FFFD;14'd9626:data <=32'h00070002;
14'd9627:data <=32'h000C0006;14'd9628:data <=32'h00120007;14'd9629:data <=32'h00170005;
14'd9630:data <=32'h001B0001;14'd9631:data <=32'h001CFFFD;14'd9632:data <=32'h001CFFFA;
14'd9633:data <=32'h001CFFF7;14'd9634:data <=32'h001CFFF6;14'd9635:data <=32'h001CFFF5;
14'd9636:data <=32'h001EFFF3;14'd9637:data <=32'h0021FFF0;14'd9638:data <=32'h0023FFEB;
14'd9639:data <=32'h0023FFE4;14'd9640:data <=32'h0021FFDC;14'd9641:data <=32'h001CFFD5;
14'd9642:data <=32'h0015FFD0;14'd9643:data <=32'h000EFFCD;14'd9644:data <=32'h0005FFCC;
14'd9645:data <=32'hFFFEFFCD;14'd9646:data <=32'hFFF7FFD0;14'd9647:data <=32'hFFF2FFD3;
14'd9648:data <=32'hFFEFFFD7;14'd9649:data <=32'hFFECFFDB;14'd9650:data <=32'hFFEAFFDF;
14'd9651:data <=32'hFFEAFFE3;14'd9652:data <=32'hFFEBFFE6;14'd9653:data <=32'hFFEEFFE8;
14'd9654:data <=32'hFFF2FFE8;14'd9655:data <=32'hFFF5FFE5;14'd9656:data <=32'hFFF7FFDE;
14'd9657:data <=32'hFFF5FFD5;14'd9658:data <=32'hFFEEFFCB;14'd9659:data <=32'hFFE2FFC4;
14'd9660:data <=32'hFFD1FFC0;14'd9661:data <=32'hFFBEFFC2;14'd9662:data <=32'hFFABFFCB;
14'd9663:data <=32'hFF9AFFDA;14'd9664:data <=32'hFFB50007;14'd9665:data <=32'hFFAE0010;
14'd9666:data <=32'hFFAE0012;14'd9667:data <=32'hFFA4FFF8;14'd9668:data <=32'hFF8C001B;
14'd9669:data <=32'hFF910030;14'd9670:data <=32'hFF9B0044;14'd9671:data <=32'hFFA90056;
14'd9672:data <=32'hFFBB0065;14'd9673:data <=32'hFFD1006E;14'd9674:data <=32'hFFE80071;
14'd9675:data <=32'hFFFE006F;14'd9676:data <=32'h00110066;14'd9677:data <=32'h0020005B;
14'd9678:data <=32'h0029004E;14'd9679:data <=32'h002F0041;14'd9680:data <=32'h00320036;
14'd9681:data <=32'h0034002D;14'd9682:data <=32'h00350025;14'd9683:data <=32'h0037001D;
14'd9684:data <=32'h00370015;14'd9685:data <=32'h0036000D;14'd9686:data <=32'h00330004;
14'd9687:data <=32'h002EFFFD;14'd9688:data <=32'h0028FFF7;14'd9689:data <=32'h0022FFF4;
14'd9690:data <=32'h001BFFF2;14'd9691:data <=32'h0016FFF2;14'd9692:data <=32'h0011FFF3;
14'd9693:data <=32'h000CFFF5;14'd9694:data <=32'h0008FFF7;14'd9695:data <=32'h0004FFFB;
14'd9696:data <=32'h00010000;14'd9697:data <=32'h00000007;14'd9698:data <=32'h0002000F;
14'd9699:data <=32'h00070017;14'd9700:data <=32'h000F001D;14'd9701:data <=32'h001B001F;
14'd9702:data <=32'h0027001D;14'd9703:data <=32'h00340017;14'd9704:data <=32'h003D000C;
14'd9705:data <=32'h0042FFFF;14'd9706:data <=32'h0043FFF0;14'd9707:data <=32'h0040FFE3;
14'd9708:data <=32'h0039FFD7;14'd9709:data <=32'h0031FFCE;14'd9710:data <=32'h0027FFC8;
14'd9711:data <=32'h001CFFC5;14'd9712:data <=32'h0013FFC3;14'd9713:data <=32'h0009FFC4;
14'd9714:data <=32'h0001FFC6;14'd9715:data <=32'hFFFAFFCB;14'd9716:data <=32'hFFF5FFD1;
14'd9717:data <=32'hFFF3FFD7;14'd9718:data <=32'hFFF4FFDC;14'd9719:data <=32'hFFF8FFDF;
14'd9720:data <=32'hFFFCFFDF;14'd9721:data <=32'h0000FFDA;14'd9722:data <=32'h0000FFD3;
14'd9723:data <=32'hFFFCFFCA;14'd9724:data <=32'hFFF4FFC1;14'd9725:data <=32'hFFE8FFBC;
14'd9726:data <=32'hFFD9FFBB;14'd9727:data <=32'hFFCAFFBE;14'd9728:data <=32'hFFE8FFB8;
14'd9729:data <=32'hFFD3FFB1;14'd9730:data <=32'hFFC5FFB6;14'd9731:data <=32'hFFCBFFDB;
14'd9732:data <=32'hFFB2FFF2;14'd9733:data <=32'hFFB2FFFD;14'd9734:data <=32'hFFB40007;
14'd9735:data <=32'hFFB70010;14'd9736:data <=32'hFFBC0018;14'd9737:data <=32'hFFC20020;
14'd9738:data <=32'hFFC90025;14'd9739:data <=32'hFFD10028;14'd9740:data <=32'hFFD60029;
14'd9741:data <=32'hFFDA0029;14'd9742:data <=32'hFFDC0029;14'd9743:data <=32'hFFDC002B;
14'd9744:data <=32'hFFDD0031;14'd9745:data <=32'hFFE00037;14'd9746:data <=32'hFFE50040;
14'd9747:data <=32'hFFEF0046;14'd9748:data <=32'hFFFB004A;14'd9749:data <=32'h0009004A;
14'd9750:data <=32'h00170046;14'd9751:data <=32'h0022003E;14'd9752:data <=32'h002B0035;
14'd9753:data <=32'h00310029;14'd9754:data <=32'h0034001E;14'd9755:data <=32'h00340012;
14'd9756:data <=32'h00320007;14'd9757:data <=32'h002CFFFD;14'd9758:data <=32'h0025FFF4;
14'd9759:data <=32'h001AFFEF;14'd9760:data <=32'h000EFFED;14'd9761:data <=32'h0003FFEF;
14'd9762:data <=32'hFFF8FFF6;14'd9763:data <=32'hFFF10000;14'd9764:data <=32'hFFEF000D;
14'd9765:data <=32'hFFF20019;14'd9766:data <=32'hFFFA0024;14'd9767:data <=32'h0005002B;
14'd9768:data <=32'h0011002E;14'd9769:data <=32'h001D002D;14'd9770:data <=32'h00280029;
14'd9771:data <=32'h00300023;14'd9772:data <=32'h0037001B;14'd9773:data <=32'h003C0013;
14'd9774:data <=32'h0040000A;14'd9775:data <=32'h00420002;14'd9776:data <=32'h0044FFF9;
14'd9777:data <=32'h0044FFEF;14'd9778:data <=32'h0043FFE5;14'd9779:data <=32'h003FFFDC;
14'd9780:data <=32'h003AFFD4;14'd9781:data <=32'h0035FFCD;14'd9782:data <=32'h002FFFC7;
14'd9783:data <=32'h002AFFC2;14'd9784:data <=32'h0024FFBC;14'd9785:data <=32'h001EFFB6;
14'd9786:data <=32'h0016FFAF;14'd9787:data <=32'h000BFFA9;14'd9788:data <=32'hFFFDFFA4;
14'd9789:data <=32'hFFEEFFA2;14'd9790:data <=32'hFFDCFFA6;14'd9791:data <=32'hFFCCFFAE;
14'd9792:data <=32'h0027FFCD;14'd9793:data <=32'h001EFFB6;14'd9794:data <=32'h0008FFA8;
14'd9795:data <=32'hFFC6FFCA;14'd9796:data <=32'hFFAFFFE6;14'd9797:data <=32'hFFB3FFF4;
14'd9798:data <=32'hFFBB0000;14'd9799:data <=32'hFFC40007;14'd9800:data <=32'hFFCD000D;
14'd9801:data <=32'hFFD6000F;14'd9802:data <=32'hFFDF000E;14'd9803:data <=32'hFFE6000B;
14'd9804:data <=32'hFFEA0004;14'd9805:data <=32'hFFE9FFFD;14'd9806:data <=32'hFFE5FFF7;
14'd9807:data <=32'hFFDDFFF4;14'd9808:data <=32'hFFD2FFF6;14'd9809:data <=32'hFFC9FFFC;
14'd9810:data <=32'hFFC20007;14'd9811:data <=32'hFFC00015;14'd9812:data <=32'hFFC30023;
14'd9813:data <=32'hFFC9002F;14'd9814:data <=32'hFFD40039;14'd9815:data <=32'hFFE0003F;
14'd9816:data <=32'hFFEC0042;14'd9817:data <=32'hFFF80042;14'd9818:data <=32'h00030040;
14'd9819:data <=32'h000E003B;14'd9820:data <=32'h00160034;14'd9821:data <=32'h001D002C;
14'd9822:data <=32'h00220021;14'd9823:data <=32'h00230017;14'd9824:data <=32'h0020000C;
14'd9825:data <=32'h001A0004;14'd9826:data <=32'h0012FFFF;14'd9827:data <=32'h000AFFFD;
14'd9828:data <=32'h0002FFFF;14'd9829:data <=32'hFFFD0003;14'd9830:data <=32'hFFFA0009;
14'd9831:data <=32'hFFF9000E;14'd9832:data <=32'hFFF90013;14'd9833:data <=32'hFFFA0017;
14'd9834:data <=32'hFFFB001A;14'd9835:data <=32'hFFFC001E;14'd9836:data <=32'hFFFD0023;
14'd9837:data <=32'h00000029;14'd9838:data <=32'h00050030;14'd9839:data <=32'h000E0037;
14'd9840:data <=32'h0019003B;14'd9841:data <=32'h0026003D;14'd9842:data <=32'h0035003B;
14'd9843:data <=32'h00440036;14'd9844:data <=32'h0051002D;14'd9845:data <=32'h005D0020;
14'd9846:data <=32'h00670011;14'd9847:data <=32'h006E0000;14'd9848:data <=32'h0072FFEC;
14'd9849:data <=32'h0072FFD6;14'd9850:data <=32'h006DFFBF;14'd9851:data <=32'h0062FFA8;
14'd9852:data <=32'h0050FF94;14'd9853:data <=32'h0039FF84;14'd9854:data <=32'h001EFF7B;
14'd9855:data <=32'h0001FF7B;14'd9856:data <=32'h0025FFDA;14'd9857:data <=32'h0027FFCB;
14'd9858:data <=32'h0022FFB4;14'd9859:data <=32'hFFF2FF8D;14'd9860:data <=32'hFFCCFFA7;
14'd9861:data <=32'hFFC3FFB7;14'd9862:data <=32'hFFBFFFC7;14'd9863:data <=32'hFFBEFFD5;
14'd9864:data <=32'hFFC0FFE2;14'd9865:data <=32'hFFC5FFED;14'd9866:data <=32'hFFCBFFF6;
14'd9867:data <=32'hFFD3FFFB;14'd9868:data <=32'hFFDBFFFD;14'd9869:data <=32'hFFE1FFFA;
14'd9870:data <=32'hFFE3FFF7;14'd9871:data <=32'hFFE2FFF3;14'd9872:data <=32'hFFDFFFF1;
14'd9873:data <=32'hFFD9FFF1;14'd9874:data <=32'hFFD3FFF5;14'd9875:data <=32'hFFD0FFFB;
14'd9876:data <=32'hFFCF0003;14'd9877:data <=32'hFFD0000B;14'd9878:data <=32'hFFD40011;
14'd9879:data <=32'hFFD80015;14'd9880:data <=32'hFFDD0017;14'd9881:data <=32'hFFE00019;
14'd9882:data <=32'hFFE3001A;14'd9883:data <=32'hFFE6001C;14'd9884:data <=32'hFFE9001D;
14'd9885:data <=32'hFFEC001F;14'd9886:data <=32'hFFF00020;14'd9887:data <=32'hFFF4001F;
14'd9888:data <=32'hFFF7001E;14'd9889:data <=32'hFFF9001C;14'd9890:data <=32'hFFFB001B;
14'd9891:data <=32'hFFFC001A;14'd9892:data <=32'hFFFD001A;14'd9893:data <=32'hFFFF001B;
14'd9894:data <=32'h0002001A;14'd9895:data <=32'h00040018;14'd9896:data <=32'h00070014;
14'd9897:data <=32'h0007000F;14'd9898:data <=32'h0004000A;14'd9899:data <=32'hFFFF0007;
14'd9900:data <=32'hFFF70006;14'd9901:data <=32'hFFEF0009;14'd9902:data <=32'hFFE70010;
14'd9903:data <=32'hFFE2001B;14'd9904:data <=32'hFFE20029;14'd9905:data <=32'hFFE60037;
14'd9906:data <=32'hFFEF0044;14'd9907:data <=32'hFFFC004F;14'd9908:data <=32'h000B0057;
14'd9909:data <=32'h001E005A;14'd9910:data <=32'h0031005A;14'd9911:data <=32'h00460055;
14'd9912:data <=32'h005A004B;14'd9913:data <=32'h006D003B;14'd9914:data <=32'h007C0026;
14'd9915:data <=32'h0085000D;14'd9916:data <=32'h0088FFF1;14'd9917:data <=32'h0083FFD5;
14'd9918:data <=32'h0076FFBC;14'd9919:data <=32'h0064FFA7;14'd9920:data <=32'h0050FFD0;
14'd9921:data <=32'h004EFFBF;14'd9922:data <=32'h004EFFB2;14'd9923:data <=32'h0057FFAC;
14'd9924:data <=32'h0033FFB1;14'd9925:data <=32'h0028FFAE;14'd9926:data <=32'h001DFFAC;
14'd9927:data <=32'h0013FFAA;14'd9928:data <=32'h0008FFAA;14'd9929:data <=32'hFFFCFFAB;
14'd9930:data <=32'hFFF2FFAE;14'd9931:data <=32'hFFE8FFB3;14'd9932:data <=32'hFFE0FFB9;
14'd9933:data <=32'hFFD9FFBE;14'd9934:data <=32'hFFD2FFC4;14'd9935:data <=32'hFFCCFFCB;
14'd9936:data <=32'hFFC5FFD3;14'd9937:data <=32'hFFBFFFDD;14'd9938:data <=32'hFFBCFFEA;
14'd9939:data <=32'hFFBBFFF8;14'd9940:data <=32'hFFC00005;14'd9941:data <=32'hFFC90010;
14'd9942:data <=32'hFFD40018;14'd9943:data <=32'hFFE0001A;14'd9944:data <=32'hFFEB0019;
14'd9945:data <=32'hFFF30014;14'd9946:data <=32'hFFF8000D;14'd9947:data <=32'hFFFA0006;
14'd9948:data <=32'hFFF90000;14'd9949:data <=32'hFFF6FFFC;14'd9950:data <=32'hFFF2FFF9;
14'd9951:data <=32'hFFEEFFF7;14'd9952:data <=32'hFFE9FFF7;14'd9953:data <=32'hFFE3FFF8;
14'd9954:data <=32'hFFDFFFFC;14'd9955:data <=32'hFFDB0001;14'd9956:data <=32'hFFD80008;
14'd9957:data <=32'hFFD8000F;14'd9958:data <=32'hFFDB0017;14'd9959:data <=32'hFFE1001D;
14'd9960:data <=32'hFFE80020;14'd9961:data <=32'hFFEF0020;14'd9962:data <=32'hFFF4001D;
14'd9963:data <=32'hFFF70018;14'd9964:data <=32'hFFF60013;14'd9965:data <=32'hFFF20010;
14'd9966:data <=32'hFFED0010;14'd9967:data <=32'hFFE70012;14'd9968:data <=32'hFFE30019;
14'd9969:data <=32'hFFE10021;14'd9970:data <=32'hFFE1002A;14'd9971:data <=32'hFFE50033;
14'd9972:data <=32'hFFEB003C;14'd9973:data <=32'hFFF30043;14'd9974:data <=32'hFFFD0049;
14'd9975:data <=32'h0008004E;14'd9976:data <=32'h00150050;14'd9977:data <=32'h00240050;
14'd9978:data <=32'h0032004C;14'd9979:data <=32'h00410044;14'd9980:data <=32'h004C0039;
14'd9981:data <=32'h0055002B;14'd9982:data <=32'h0059001C;14'd9983:data <=32'h0059000E;
14'd9984:data <=32'h0079001B;14'd9985:data <=32'h00840004;14'd9986:data <=32'h0082FFF4;
14'd9987:data <=32'h005A0011;14'd9988:data <=32'h00480015;14'd9989:data <=32'h0050000E;
14'd9990:data <=32'h00580003;14'd9991:data <=32'h005FFFF5;14'd9992:data <=32'h0060FFE4;
14'd9993:data <=32'h005EFFD2;14'd9994:data <=32'h0057FFC1;14'd9995:data <=32'h004CFFB2;
14'd9996:data <=32'h003EFFA5;14'd9997:data <=32'h002EFF9A;14'd9998:data <=32'h001CFF93;
14'd9999:data <=32'h0007FF90;14'd10000:data <=32'hFFF1FF91;14'd10001:data <=32'hFFDBFF98;
14'd10002:data <=32'hFFC7FFA6;14'd10003:data <=32'hFFB8FFB8;14'd10004:data <=32'hFFB0FFCE;
14'd10005:data <=32'hFFAFFFE4;14'd10006:data <=32'hFFB4FFF8;14'd10007:data <=32'hFFBF0008;
14'd10008:data <=32'hFFCC0013;14'd10009:data <=32'hFFDA0019;14'd10010:data <=32'hFFE80019;
14'd10011:data <=32'hFFF30016;14'd10012:data <=32'hFFFB0011;14'd10013:data <=32'h0002000B;
14'd10014:data <=32'h00060003;14'd10015:data <=32'h0008FFFC;14'd10016:data <=32'h0007FFF3;
14'd10017:data <=32'h0004FFEB;14'd10018:data <=32'hFFFFFFE5;14'd10019:data <=32'hFFF7FFE1;
14'd10020:data <=32'hFFEFFFDF;14'd10021:data <=32'hFFE6FFE0;14'd10022:data <=32'hFFDEFFE4;
14'd10023:data <=32'hFFD9FFE9;14'd10024:data <=32'hFFD5FFEF;14'd10025:data <=32'hFFD3FFF4;
14'd10026:data <=32'hFFD1FFF9;14'd10027:data <=32'hFFCFFFFC;14'd10028:data <=32'hFFCD0000;
14'd10029:data <=32'hFFC90005;14'd10030:data <=32'hFFC6000C;14'd10031:data <=32'hFFC30015;
14'd10032:data <=32'hFFC30020;14'd10033:data <=32'hFFC6002B;14'd10034:data <=32'hFFCD0036;
14'd10035:data <=32'hFFD6003F;14'd10036:data <=32'hFFE20044;14'd10037:data <=32'hFFED0047;
14'd10038:data <=32'hFFF80048;14'd10039:data <=32'h00020046;14'd10040:data <=32'h000B0043;
14'd10041:data <=32'h0012003F;14'd10042:data <=32'h00190039;14'd10043:data <=32'h001E0034;
14'd10044:data <=32'h0021002D;14'd10045:data <=32'h00220026;14'd10046:data <=32'h00210021;
14'd10047:data <=32'h001E001D;14'd10048:data <=32'h0034005F;14'd10049:data <=32'h004A005A;
14'd10050:data <=32'h00540049;14'd10051:data <=32'h00220026;14'd10052:data <=32'h000E0037;
14'd10053:data <=32'h001A003E;14'd10054:data <=32'h00290041;14'd10055:data <=32'h003B003E;
14'd10056:data <=32'h004B0036;14'd10057:data <=32'h00580029;14'd10058:data <=32'h0062001A;
14'd10059:data <=32'h00680008;14'd10060:data <=32'h006AFFF5;14'd10061:data <=32'h0068FFE1;
14'd10062:data <=32'h0062FFCE;14'd10063:data <=32'h0057FFBB;14'd10064:data <=32'h0048FFAC;
14'd10065:data <=32'h0034FFA1;14'd10066:data <=32'h001EFF9C;14'd10067:data <=32'h0008FF9E;
14'd10068:data <=32'hFFF5FFA5;14'd10069:data <=32'hFFE5FFB1;14'd10070:data <=32'hFFDBFFBF;
14'd10071:data <=32'hFFD5FFCD;14'd10072:data <=32'hFFD5FFDA;14'd10073:data <=32'hFFD6FFE5;
14'd10074:data <=32'hFFD9FFEE;14'd10075:data <=32'hFFDDFFF6;14'd10076:data <=32'hFFE1FFFB;
14'd10077:data <=32'hFFE60001;14'd10078:data <=32'hFFEC0005;14'd10079:data <=32'hFFF30008;
14'd10080:data <=32'hFFFA0008;14'd10081:data <=32'h00020006;14'd10082:data <=32'h00090001;
14'd10083:data <=32'h000DFFFB;14'd10084:data <=32'h000FFFF4;14'd10085:data <=32'h0010FFEC;
14'd10086:data <=32'h000EFFE4;14'd10087:data <=32'h000BFFDD;14'd10088:data <=32'h0006FFD6;
14'd10089:data <=32'h0000FFCF;14'd10090:data <=32'hFFF7FFC9;14'd10091:data <=32'hFFECFFC4;
14'd10092:data <=32'hFFDFFFC0;14'd10093:data <=32'hFFCFFFC2;14'd10094:data <=32'hFFBEFFC7;
14'd10095:data <=32'hFFAEFFD2;14'd10096:data <=32'hFFA1FFE2;14'd10097:data <=32'hFF99FFF6;
14'd10098:data <=32'hFF97000C;14'd10099:data <=32'hFF9C0021;14'd10100:data <=32'hFFA50034;
14'd10101:data <=32'hFFB30042;14'd10102:data <=32'hFFC3004D;14'd10103:data <=32'hFFD30053;
14'd10104:data <=32'hFFE30055;14'd10105:data <=32'hFFF20054;14'd10106:data <=32'h0000004F;
14'd10107:data <=32'h000C0048;14'd10108:data <=32'h0014003F;14'd10109:data <=32'h00190034;
14'd10110:data <=32'h001A0029;14'd10111:data <=32'h00160021;14'd10112:data <=32'hFFF6003A;
14'd10113:data <=32'hFFFB0042;14'd10114:data <=32'h00080045;14'd10115:data <=32'h001C002C;
14'd10116:data <=32'h00040037;14'd10117:data <=32'h000A003C;14'd10118:data <=32'h00130040;
14'd10119:data <=32'h001F0040;14'd10120:data <=32'h002A003D;14'd10121:data <=32'h00340037;
14'd10122:data <=32'h003C002F;14'd10123:data <=32'h00410025;14'd10124:data <=32'h0045001C;
14'd10125:data <=32'h00480012;14'd10126:data <=32'h004A0008;14'd10127:data <=32'h0049FFFD;
14'd10128:data <=32'h0046FFF2;14'd10129:data <=32'h0041FFE8;14'd10130:data <=32'h003AFFDF;
14'd10131:data <=32'h0031FFDA;14'd10132:data <=32'h0027FFD8;14'd10133:data <=32'h0020FFD8;
14'd10134:data <=32'h001AFFD9;14'd10135:data <=32'h0017FFDA;14'd10136:data <=32'h0015FFDB;
14'd10137:data <=32'h0013FFDA;14'd10138:data <=32'h000FFFD7;14'd10139:data <=32'h000AFFD5;
14'd10140:data <=32'h0003FFD4;14'd10141:data <=32'hFFFBFFD6;14'd10142:data <=32'hFFF4FFDB;
14'd10143:data <=32'hFFEFFFE1;14'd10144:data <=32'hFFECFFE9;14'd10145:data <=32'hFFEDFFF2;
14'd10146:data <=32'hFFF0FFF9;14'd10147:data <=32'hFFF6FFFF;14'd10148:data <=32'hFFFC0002;
14'd10149:data <=32'h00030003;14'd10150:data <=32'h000B0002;14'd10151:data <=32'h0013FFFF;
14'd10152:data <=32'h001BFFF9;14'd10153:data <=32'h0020FFEF;14'd10154:data <=32'h0024FFE3;
14'd10155:data <=32'h0024FFD5;14'd10156:data <=32'h001EFFC6;14'd10157:data <=32'h0013FFB8;
14'd10158:data <=32'h0004FFAD;14'd10159:data <=32'hFFF0FFA8;14'd10160:data <=32'hFFDCFFA8;
14'd10161:data <=32'hFFC8FFAE;14'd10162:data <=32'hFFB7FFBA;14'd10163:data <=32'hFFAAFFCA;
14'd10164:data <=32'hFFA2FFDB;14'd10165:data <=32'hFF9EFFEC;14'd10166:data <=32'hFF9EFFFC;
14'd10167:data <=32'hFFA1000B;14'd10168:data <=32'hFFA60018;14'd10169:data <=32'hFFAC0024;
14'd10170:data <=32'hFFB4002F;14'd10171:data <=32'hFFBD0037;14'd10172:data <=32'hFFC8003D;
14'd10173:data <=32'hFFD20041;14'd10174:data <=32'hFFDC0041;14'd10175:data <=32'hFFE30041;
14'd10176:data <=32'hFFFE0024;14'd10177:data <=32'hFFF90022;14'd10178:data <=32'hFFF40029;
14'd10179:data <=32'hFFEB0054;14'd10180:data <=32'hFFDE0062;14'd10181:data <=32'hFFEE0068;
14'd10182:data <=32'h0002006A;14'd10183:data <=32'h00160067;14'd10184:data <=32'h0028005F;
14'd10185:data <=32'h00370052;14'd10186:data <=32'h00410042;14'd10187:data <=32'h00460031;
14'd10188:data <=32'h00470021;14'd10189:data <=32'h00440014;14'd10190:data <=32'h003F0009;
14'd10191:data <=32'h00380000;14'd10192:data <=32'h0031FFF9;14'd10193:data <=32'h0029FFF5;
14'd10194:data <=32'h0020FFF3;14'd10195:data <=32'h0018FFF4;14'd10196:data <=32'h0012FFF9;
14'd10197:data <=32'h000FFFFF;14'd10198:data <=32'h000F0005;14'd10199:data <=32'h0014000B;
14'd10200:data <=32'h001A000D;14'd10201:data <=32'h0023000B;14'd10202:data <=32'h00290006;
14'd10203:data <=32'h002DFFFE;14'd10204:data <=32'h002EFFF4;14'd10205:data <=32'h002BFFEC;
14'd10206:data <=32'h0025FFE4;14'd10207:data <=32'h001DFFE0;14'd10208:data <=32'h0016FFDF;
14'd10209:data <=32'h000FFFE0;14'd10210:data <=32'h000AFFE2;14'd10211:data <=32'h0006FFE6;
14'd10212:data <=32'h0003FFEA;14'd10213:data <=32'h0003FFEE;14'd10214:data <=32'h0003FFF2;
14'd10215:data <=32'h0005FFF6;14'd10216:data <=32'h0009FFFA;14'd10217:data <=32'h000FFFFB;
14'd10218:data <=32'h0016FFF9;14'd10219:data <=32'h001CFFF4;14'd10220:data <=32'h0021FFED;
14'd10221:data <=32'h0023FFE3;14'd10222:data <=32'h0021FFD9;14'd10223:data <=32'h001CFFCF;
14'd10224:data <=32'h0014FFC7;14'd10225:data <=32'h000BFFC2;14'd10226:data <=32'h0002FFBF;
14'd10227:data <=32'hFFF9FFBF;14'd10228:data <=32'hFFF2FFC0;14'd10229:data <=32'hFFEBFFC0;
14'd10230:data <=32'hFFE4FFC0;14'd10231:data <=32'hFFDCFFC0;14'd10232:data <=32'hFFD3FFC0;
14'd10233:data <=32'hFFC8FFC2;14'd10234:data <=32'hFFBDFFC7;14'd10235:data <=32'hFFB2FFCF;
14'd10236:data <=32'hFFA7FFD9;14'd10237:data <=32'hFF9FFFE5;14'd10238:data <=32'hFF99FFF4;
14'd10239:data <=32'hFF940003;14'd10240:data <=32'hFFDD0028;14'd10241:data <=32'hFFDE0024;
14'd10242:data <=32'hFFD4001E;14'd10243:data <=32'hFF94001F;14'd10244:data <=32'hFF7F003E;
14'd10245:data <=32'hFF8E0058;14'd10246:data <=32'hFFA3006D;14'd10247:data <=32'hFFBD007C;
14'd10248:data <=32'hFFDA0083;14'd10249:data <=32'hFFF70081;14'd10250:data <=32'h00100078;
14'd10251:data <=32'h0025006B;14'd10252:data <=32'h0034005A;14'd10253:data <=32'h003D0047;
14'd10254:data <=32'h00420036;14'd10255:data <=32'h00420025;14'd10256:data <=32'h003F0016;
14'd10257:data <=32'h00390008;14'd10258:data <=32'h0030FFFE;14'd10259:data <=32'h0025FFF7;
14'd10260:data <=32'h0019FFF5;14'd10261:data <=32'h000FFFF8;14'd10262:data <=32'h0007FFFD;
14'd10263:data <=32'h00040005;14'd10264:data <=32'h0004000D;14'd10265:data <=32'h00080012;
14'd10266:data <=32'h000D0016;14'd10267:data <=32'h00130016;14'd10268:data <=32'h00180013;
14'd10269:data <=32'h001B0010;14'd10270:data <=32'h001C000D;14'd10271:data <=32'h001D000A;
14'd10272:data <=32'h001D0009;14'd10273:data <=32'h001E0008;14'd10274:data <=32'h00200006;
14'd10275:data <=32'h00220004;14'd10276:data <=32'h00240001;14'd10277:data <=32'h0025FFFE;
14'd10278:data <=32'h0025FFFA;14'd10279:data <=32'h0025FFF6;14'd10280:data <=32'h0023FFF2;
14'd10281:data <=32'h0022FFEF;14'd10282:data <=32'h0021FFEC;14'd10283:data <=32'h0020FFE9;
14'd10284:data <=32'h001EFFE6;14'd10285:data <=32'h001CFFE3;14'd10286:data <=32'h0018FFE0;
14'd10287:data <=32'h0014FFDE;14'd10288:data <=32'h000FFFDE;14'd10289:data <=32'h000BFFE0;
14'd10290:data <=32'h0009FFE3;14'd10291:data <=32'h000AFFE7;14'd10292:data <=32'h000EFFE9;
14'd10293:data <=32'h0014FFE8;14'd10294:data <=32'h001AFFE3;14'd10295:data <=32'h001FFFDA;
14'd10296:data <=32'h0020FFCE;14'd10297:data <=32'h001CFFC0;14'd10298:data <=32'h0014FFB3;
14'd10299:data <=32'h0007FFA7;14'd10300:data <=32'hFFF6FF9F;14'd10301:data <=32'hFFE3FF9B;
14'd10302:data <=32'hFFCFFF9B;14'd10303:data <=32'hFFBAFFA0;14'd10304:data <=32'hFFC7FFDF;
14'd10305:data <=32'hFFBDFFDD;14'd10306:data <=32'hFFB8FFD8;14'd10307:data <=32'hFFABFFB7;
14'd10308:data <=32'hFF83FFD0;14'd10309:data <=32'hFF7BFFEB;14'd10310:data <=32'hFF7B0006;
14'd10311:data <=32'hFF820020;14'd10312:data <=32'hFF8F0036;14'd10313:data <=32'hFFA00047;
14'd10314:data <=32'hFFB40051;14'd10315:data <=32'hFFC60056;14'd10316:data <=32'hFFD70058;
14'd10317:data <=32'hFFE60057;14'd10318:data <=32'hFFF30054;14'd10319:data <=32'hFFFF0050;
14'd10320:data <=32'h000A0049;14'd10321:data <=32'h00140042;14'd10322:data <=32'h001A0039;
14'd10323:data <=32'h001E002F;14'd10324:data <=32'h001F0026;14'd10325:data <=32'h001E001F;
14'd10326:data <=32'h001C0019;14'd10327:data <=32'h001B0015;14'd10328:data <=32'h001A0012;
14'd10329:data <=32'h0019000F;14'd10330:data <=32'h0018000C;14'd10331:data <=32'h00170008;
14'd10332:data <=32'h00130004;14'd10333:data <=32'h000E0001;14'd10334:data <=32'h00070000;
14'd10335:data <=32'h00010003;14'd10336:data <=32'hFFFC0008;14'd10337:data <=32'hFFF90010;
14'd10338:data <=32'hFFFB0019;14'd10339:data <=32'hFFFF0021;14'd10340:data <=32'h00070027;
14'd10341:data <=32'h0011002A;14'd10342:data <=32'h001A002A;14'd10343:data <=32'h00240027;
14'd10344:data <=32'h002C0022;14'd10345:data <=32'h0034001B;14'd10346:data <=32'h00390013;
14'd10347:data <=32'h003D0009;14'd10348:data <=32'h003EFFFF;14'd10349:data <=32'h003DFFF4;
14'd10350:data <=32'h0039FFEA;14'd10351:data <=32'h0031FFE1;14'd10352:data <=32'h0028FFDD;
14'd10353:data <=32'h001FFFDB;14'd10354:data <=32'h0016FFDE;14'd10355:data <=32'h0011FFE3;
14'd10356:data <=32'h000FFFE9;14'd10357:data <=32'h0012FFEF;14'd10358:data <=32'h0018FFF2;
14'd10359:data <=32'h0020FFF1;14'd10360:data <=32'h0027FFEB;14'd10361:data <=32'h002CFFE2;
14'd10362:data <=32'h002EFFD6;14'd10363:data <=32'h002CFFC9;14'd10364:data <=32'h0026FFBE;
14'd10365:data <=32'h001DFFB2;14'd10366:data <=32'h0012FFA9;14'd10367:data <=32'h0003FFA2;
14'd10368:data <=32'h0019FFAF;14'd10369:data <=32'h000AFF9B;14'd10370:data <=32'hFFFBFF94;
14'd10371:data <=32'hFFF4FFAF;14'd10372:data <=32'hFFCCFFB7;14'd10373:data <=32'hFFC2FFC2;
14'd10374:data <=32'hFFBBFFCE;14'd10375:data <=32'hFFB8FFDB;14'd10376:data <=32'hFFB8FFE6;
14'd10377:data <=32'hFFBAFFEF;14'd10378:data <=32'hFFBDFFF5;14'd10379:data <=32'hFFBEFFF9;
14'd10380:data <=32'hFFBEFFFD;14'd10381:data <=32'hFFBD0003;14'd10382:data <=32'hFFBB0009;
14'd10383:data <=32'hFFBA0012;14'd10384:data <=32'hFFBC001D;14'd10385:data <=32'hFFC00027;
14'd10386:data <=32'hFFC60030;14'd10387:data <=32'hFFCF0038;14'd10388:data <=32'hFFD8003D;
14'd10389:data <=32'hFFE30041;14'd10390:data <=32'hFFEE0044;14'd10391:data <=32'hFFF90045;
14'd10392:data <=32'h00050042;14'd10393:data <=32'h0011003D;14'd10394:data <=32'h001C0034;
14'd10395:data <=32'h00240028;14'd10396:data <=32'h0028001B;14'd10397:data <=32'h0027000C;
14'd10398:data <=32'h00200000;14'd10399:data <=32'h0016FFF7;14'd10400:data <=32'h0009FFF3;
14'd10401:data <=32'hFFFCFFF4;14'd10402:data <=32'hFFF2FFFA;14'd10403:data <=32'hFFEB0003;
14'd10404:data <=32'hFFE7000D;14'd10405:data <=32'hFFE70018;14'd10406:data <=32'hFFEA0022;
14'd10407:data <=32'hFFF0002A;14'd10408:data <=32'hFFF70031;14'd10409:data <=32'h00000036;
14'd10410:data <=32'h000A0039;14'd10411:data <=32'h0015003A;14'd10412:data <=32'h00200038;
14'd10413:data <=32'h002A0033;14'd10414:data <=32'h0033002C;14'd10415:data <=32'h00390023;
14'd10416:data <=32'h003D001A;14'd10417:data <=32'h003E0011;14'd10418:data <=32'h003D000A;
14'd10419:data <=32'h003C0005;14'd10420:data <=32'h003C0001;14'd10421:data <=32'h003DFFFD;
14'd10422:data <=32'h0041FFF8;14'd10423:data <=32'h0044FFF2;14'd10424:data <=32'h0046FFE8;
14'd10425:data <=32'h0046FFDD;14'd10426:data <=32'h0042FFD0;14'd10427:data <=32'h003BFFC5;
14'd10428:data <=32'h0032FFBB;14'd10429:data <=32'h0026FFB5;14'd10430:data <=32'h001AFFB1;
14'd10431:data <=32'h000FFFAF;14'd10432:data <=32'h0051FFE8;14'd10433:data <=32'h0056FFCB;
14'd10434:data <=32'h004AFFB2;14'd10435:data <=32'h0001FFB7;14'd10436:data <=32'hFFDEFFC2;
14'd10437:data <=32'hFFD9FFCD;14'd10438:data <=32'hFFD9FFD9;14'd10439:data <=32'hFFDBFFE3;
14'd10440:data <=32'hFFE1FFEB;14'd10441:data <=32'hFFE9FFED;14'd10442:data <=32'hFFF0FFEB;
14'd10443:data <=32'hFFF5FFE5;14'd10444:data <=32'hFFF4FFDD;14'd10445:data <=32'hFFEFFFD5;
14'd10446:data <=32'hFFE6FFD1;14'd10447:data <=32'hFFDAFFD0;14'd10448:data <=32'hFFCDFFD3;
14'd10449:data <=32'hFFC3FFDA;14'd10450:data <=32'hFFBBFFE5;14'd10451:data <=32'hFFB5FFF0;
14'd10452:data <=32'hFFB2FFFD;14'd10453:data <=32'hFFB2000B;14'd10454:data <=32'hFFB50019;
14'd10455:data <=32'hFFBB0027;14'd10456:data <=32'hFFC50033;14'd10457:data <=32'hFFD2003C;
14'd10458:data <=32'hFFE20040;14'd10459:data <=32'hFFF20041;14'd10460:data <=32'h0001003C;
14'd10461:data <=32'h000C0032;14'd10462:data <=32'h00130026;14'd10463:data <=32'h0016001A;
14'd10464:data <=32'h0014000F;14'd10465:data <=32'h000F0007;14'd10466:data <=32'h00080002;
14'd10467:data <=32'h0002FFFF;14'd10468:data <=32'hFFFCFFFE;14'd10469:data <=32'hFFF7FFFF;
14'd10470:data <=32'hFFF20001;14'd10471:data <=32'hFFED0004;14'd10472:data <=32'hFFE80007;
14'd10473:data <=32'hFFE4000C;14'd10474:data <=32'hFFE10013;14'd10475:data <=32'hFFE0001C;
14'd10476:data <=32'hFFE00025;14'd10477:data <=32'hFFE3002E;14'd10478:data <=32'hFFE80037;
14'd10479:data <=32'hFFF0003F;14'd10480:data <=32'hFFF90046;14'd10481:data <=32'h0003004B;
14'd10482:data <=32'h000E004F;14'd10483:data <=32'h001B0052;14'd10484:data <=32'h002A0053;
14'd10485:data <=32'h003B0051;14'd10486:data <=32'h004D004A;14'd10487:data <=32'h005E003F;
14'd10488:data <=32'h006E002E;14'd10489:data <=32'h00790018;14'd10490:data <=32'h007EFFFF;
14'd10491:data <=32'h007BFFE5;14'd10492:data <=32'h0073FFCE;14'd10493:data <=32'h0064FFBA;
14'd10494:data <=32'h0052FFAB;14'd10495:data <=32'h003FFFA2;14'd10496:data <=32'h003C0009;
14'd10497:data <=32'h004CFFFA;14'd10498:data <=32'h0056FFDF;14'd10499:data <=32'h0032FFA2;
14'd10500:data <=32'h0006FFA6;14'd10501:data <=32'hFFF7FFB0;14'd10502:data <=32'hFFEDFFBC;
14'd10503:data <=32'hFFE7FFC9;14'd10504:data <=32'hFFE7FFD6;14'd10505:data <=32'hFFEBFFE0;
14'd10506:data <=32'hFFF1FFE5;14'd10507:data <=32'hFFF9FFE6;14'd10508:data <=32'hFFFDFFE2;
14'd10509:data <=32'hFFFEFFDD;14'd10510:data <=32'hFFFCFFD7;14'd10511:data <=32'hFFF6FFD2;
14'd10512:data <=32'hFFEFFFD1;14'd10513:data <=32'hFFE8FFD2;14'd10514:data <=32'hFFE1FFD4;
14'd10515:data <=32'hFFDBFFD8;14'd10516:data <=32'hFFD6FFDC;14'd10517:data <=32'hFFD1FFE2;
14'd10518:data <=32'hFFCDFFE8;14'd10519:data <=32'hFFCAFFF0;14'd10520:data <=32'hFFC9FFF9;
14'd10521:data <=32'hFFCA0002;14'd10522:data <=32'hFFCD000A;14'd10523:data <=32'hFFD30011;
14'd10524:data <=32'hFFDA0015;14'd10525:data <=32'hFFE10016;14'd10526:data <=32'hFFE60016;
14'd10527:data <=32'hFFEA0014;14'd10528:data <=32'hFFEC0013;14'd10529:data <=32'hFFED0012;
14'd10530:data <=32'hFFEE0013;14'd10531:data <=32'hFFF00014;14'd10532:data <=32'hFFF40015;
14'd10533:data <=32'hFFF80014;14'd10534:data <=32'hFFFC0011;14'd10535:data <=32'hFFFE000C;
14'd10536:data <=32'hFFFE0006;14'd10537:data <=32'hFFFBFFFF;14'd10538:data <=32'hFFF6FFFA;
14'd10539:data <=32'hFFEEFFF8;14'd10540:data <=32'hFFE5FFF8;14'd10541:data <=32'hFFDBFFFB;
14'd10542:data <=32'hFFD30002;14'd10543:data <=32'hFFCC000C;14'd10544:data <=32'hFFC60017;
14'd10545:data <=32'hFFC30025;14'd10546:data <=32'hFFC40035;14'd10547:data <=32'hFFC80046;
14'd10548:data <=32'hFFD20058;14'd10549:data <=32'hFFE10069;14'd10550:data <=32'hFFF60075;
14'd10551:data <=32'h000F007C;14'd10552:data <=32'h002B007C;14'd10553:data <=32'h00460073;
14'd10554:data <=32'h005E0063;14'd10555:data <=32'h0071004D;14'd10556:data <=32'h007C0035;
14'd10557:data <=32'h0081001B;14'd10558:data <=32'h007F0003;14'd10559:data <=32'h0079FFED;
14'd10560:data <=32'h004F000C;14'd10561:data <=32'h005A0001;14'd10562:data <=32'h0067FFF6;
14'd10563:data <=32'h0079FFE8;14'd10564:data <=32'h0056FFDA;14'd10565:data <=32'h004CFFD1;
14'd10566:data <=32'h0042FFCB;14'd10567:data <=32'h0038FFC7;14'd10568:data <=32'h002FFFC5;
14'd10569:data <=32'h0028FFC4;14'd10570:data <=32'h0023FFC3;14'd10571:data <=32'h001EFFC0;
14'd10572:data <=32'h0017FFBC;14'd10573:data <=32'h000FFFB8;14'd10574:data <=32'h0004FFB6;
14'd10575:data <=32'hFFF8FFB7;14'd10576:data <=32'hFFECFFBC;14'd10577:data <=32'hFFE2FFC4;
14'd10578:data <=32'hFFDAFFCE;14'd10579:data <=32'hFFD7FFD9;14'd10580:data <=32'hFFD7FFE3;
14'd10581:data <=32'hFFDAFFEB;14'd10582:data <=32'hFFDDFFF2;14'd10583:data <=32'hFFE1FFF6;
14'd10584:data <=32'hFFE5FFF9;14'd10585:data <=32'hFFEAFFFB;14'd10586:data <=32'hFFEEFFFC;
14'd10587:data <=32'hFFF2FFFB;14'd10588:data <=32'hFFF6FFF8;14'd10589:data <=32'hFFF7FFF4;
14'd10590:data <=32'hFFF6FFEE;14'd10591:data <=32'hFFF3FFEA;14'd10592:data <=32'hFFEDFFE8;
14'd10593:data <=32'hFFE6FFE8;14'd10594:data <=32'hFFDFFFEC;14'd10595:data <=32'hFFDAFFF2;
14'd10596:data <=32'hFFD8FFFA;14'd10597:data <=32'hFFD90002;14'd10598:data <=32'hFFDD0008;
14'd10599:data <=32'hFFE3000B;14'd10600:data <=32'hFFE9000C;14'd10601:data <=32'hFFEE0009;
14'd10602:data <=32'hFFF00005;14'd10603:data <=32'hFFF00001;14'd10604:data <=32'hFFEEFFFC;
14'd10605:data <=32'hFFE9FFF9;14'd10606:data <=32'hFFE4FFF8;14'd10607:data <=32'hFFDDFFF8;
14'd10608:data <=32'hFFD6FFFA;14'd10609:data <=32'hFFCEFFFF;14'd10610:data <=32'hFFC70007;
14'd10611:data <=32'hFFC00011;14'd10612:data <=32'hFFBC001F;14'd10613:data <=32'hFFBD002F;
14'd10614:data <=32'hFFC1003F;14'd10615:data <=32'hFFCC004F;14'd10616:data <=32'hFFDA005B;
14'd10617:data <=32'hFFEC0063;14'd10618:data <=32'hFFFF0066;14'd10619:data <=32'h00100063;
14'd10620:data <=32'h001F005D;14'd10621:data <=32'h002C0056;14'd10622:data <=32'h0035004E;
14'd10623:data <=32'h003E0045;14'd10624:data <=32'h00520052;14'd10625:data <=32'h00650047;
14'd10626:data <=32'h006E003D;14'd10627:data <=32'h004A004B;14'd10628:data <=32'h003B0044;
14'd10629:data <=32'h0046003E;14'd10630:data <=32'h00510035;14'd10631:data <=32'h005B002B;
14'd10632:data <=32'h0062001E;14'd10633:data <=32'h0069000F;14'd10634:data <=32'h006EFFFE;
14'd10635:data <=32'h0070FFEA;14'd10636:data <=32'h006CFFD5;14'd10637:data <=32'h0063FFC0;
14'd10638:data <=32'h0053FFAD;14'd10639:data <=32'h003FFF9F;14'd10640:data <=32'h0027FF98;
14'd10641:data <=32'h000FFF99;14'd10642:data <=32'hFFF9FFA0;14'd10643:data <=32'hFFE8FFAB;
14'd10644:data <=32'hFFDBFFBA;14'd10645:data <=32'hFFD4FFCA;14'd10646:data <=32'hFFD1FFD9;
14'd10647:data <=32'hFFD2FFE7;14'd10648:data <=32'hFFD7FFF4;14'd10649:data <=32'hFFDDFFFE;
14'd10650:data <=32'hFFE60006;14'd10651:data <=32'hFFF0000A;14'd10652:data <=32'hFFFB000B;
14'd10653:data <=32'h00050007;14'd10654:data <=32'h000D0000;14'd10655:data <=32'h0012FFF7;
14'd10656:data <=32'h0012FFEC;14'd10657:data <=32'h000FFFE4;14'd10658:data <=32'h0008FFDD;
14'd10659:data <=32'h0000FFDA;14'd10660:data <=32'hFFF9FFD9;14'd10661:data <=32'hFFF3FFDA;
14'd10662:data <=32'hFFEFFFDD;14'd10663:data <=32'hFFECFFDF;14'd10664:data <=32'hFFE9FFE0;
14'd10665:data <=32'hFFE6FFE0;14'd10666:data <=32'hFFE3FFE0;14'd10667:data <=32'hFFDEFFE1;
14'd10668:data <=32'hFFD8FFE3;14'd10669:data <=32'hFFD2FFE6;14'd10670:data <=32'hFFCDFFEC;
14'd10671:data <=32'hFFCAFFF2;14'd10672:data <=32'hFFC7FFF9;14'd10673:data <=32'hFFC5FFFF;
14'd10674:data <=32'hFFC50006;14'd10675:data <=32'hFFC4000E;14'd10676:data <=32'hFFC50015;
14'd10677:data <=32'hFFC7001E;14'd10678:data <=32'hFFCB0026;14'd10679:data <=32'hFFD1002D;
14'd10680:data <=32'hFFD90033;14'd10681:data <=32'hFFE10035;14'd10682:data <=32'hFFEA0035;
14'd10683:data <=32'hFFF00032;14'd10684:data <=32'hFFF3002F;14'd10685:data <=32'hFFF4002C;
14'd10686:data <=32'hFFF1002C;14'd10687:data <=32'hFFEF002F;14'd10688:data <=32'hFFF70070;
14'd10689:data <=32'h000C0078;14'd10690:data <=32'h001C0071;14'd10691:data <=32'hFFF90042;
14'd10692:data <=32'hFFE5004A;14'd10693:data <=32'hFFF00055;14'd10694:data <=32'hFFFF005D;
14'd10695:data <=32'h000F0062;14'd10696:data <=32'h00220064;14'd10697:data <=32'h00360061;
14'd10698:data <=32'h004A0059;14'd10699:data <=32'h005E004C;14'd10700:data <=32'h006E0038;
14'd10701:data <=32'h00780020;14'd10702:data <=32'h007B0006;14'd10703:data <=32'h0077FFEC;
14'd10704:data <=32'h006BFFD5;14'd10705:data <=32'h005AFFC4;14'd10706:data <=32'h0048FFB9;
14'd10707:data <=32'h0034FFB3;14'd10708:data <=32'h0022FFB3;14'd10709:data <=32'h0012FFB6;
14'd10710:data <=32'h0005FFBB;14'd10711:data <=32'hFFFAFFC2;14'd10712:data <=32'hFFF1FFCB;
14'd10713:data <=32'hFFEAFFD5;14'd10714:data <=32'hFFE7FFE0;14'd10715:data <=32'hFFE6FFEB;
14'd10716:data <=32'hFFE9FFF5;14'd10717:data <=32'hFFEFFFFD;14'd10718:data <=32'hFFF60002;
14'd10719:data <=32'hFFFE0005;14'd10720:data <=32'h00050004;14'd10721:data <=32'h000B0002;
14'd10722:data <=32'h000FFFFE;14'd10723:data <=32'h0013FFFB;14'd10724:data <=32'h0016FFF8;
14'd10725:data <=32'h0019FFF3;14'd10726:data <=32'h001CFFEE;14'd10727:data <=32'h001FFFE6;
14'd10728:data <=32'h0020FFDD;14'd10729:data <=32'h001EFFD2;14'd10730:data <=32'h0018FFC6;
14'd10731:data <=32'h000FFFBB;14'd10732:data <=32'h0001FFB4;14'd10733:data <=32'hFFF1FFB0;
14'd10734:data <=32'hFFDFFFB0;14'd10735:data <=32'hFFD0FFB6;14'd10736:data <=32'hFFC1FFBF;
14'd10737:data <=32'hFFB6FFCB;14'd10738:data <=32'hFFADFFD9;14'd10739:data <=32'hFFA8FFE8;
14'd10740:data <=32'hFFA7FFF8;14'd10741:data <=32'hFFA90008;14'd10742:data <=32'hFFAD0017;
14'd10743:data <=32'hFFB60023;14'd10744:data <=32'hFFC2002D;14'd10745:data <=32'hFFD00033;
14'd10746:data <=32'hFFDE0033;14'd10747:data <=32'hFFE9002F;14'd10748:data <=32'hFFF10027;
14'd10749:data <=32'hFFF4001E;14'd10750:data <=32'hFFF10016;14'd10751:data <=32'hFFEA0012;
14'd10752:data <=32'hFFC70027;14'd10753:data <=32'hFFC60034;14'd10754:data <=32'hFFD2003F;
14'd10755:data <=32'hFFED002B;14'd10756:data <=32'hFFD4002E;14'd10757:data <=32'hFFD70037;
14'd10758:data <=32'hFFDD0040;14'd10759:data <=32'hFFE60047;14'd10760:data <=32'hFFEF004E;
14'd10761:data <=32'hFFFB0053;14'd10762:data <=32'h00080057;14'd10763:data <=32'h00180056;
14'd10764:data <=32'h00270051;14'd10765:data <=32'h00360048;14'd10766:data <=32'h0041003C;
14'd10767:data <=32'h0047002D;14'd10768:data <=32'h0049001F;14'd10769:data <=32'h00470012;
14'd10770:data <=32'h00430008;14'd10771:data <=32'h003E0000;14'd10772:data <=32'h003AFFFB;
14'd10773:data <=32'h0037FFF6;14'd10774:data <=32'h0034FFF2;14'd10775:data <=32'h0031FFEC;
14'd10776:data <=32'h002DFFE6;14'd10777:data <=32'h0027FFE2;14'd10778:data <=32'h0020FFDE;
14'd10779:data <=32'h0019FFDD;14'd10780:data <=32'h0012FFDD;14'd10781:data <=32'h000BFFDF;
14'd10782:data <=32'h0005FFE2;14'd10783:data <=32'h0001FFE6;14'd10784:data <=32'hFFFDFFEB;
14'd10785:data <=32'hFFFBFFF0;14'd10786:data <=32'hFFFAFFF6;14'd10787:data <=32'hFFFAFFFD;
14'd10788:data <=32'hFFFD0005;14'd10789:data <=32'h0003000C;14'd10790:data <=32'h000D0010;
14'd10791:data <=32'h001A0012;14'd10792:data <=32'h0027000E;14'd10793:data <=32'h00330005;
14'd10794:data <=32'h003CFFF7;14'd10795:data <=32'h0040FFE6;14'd10796:data <=32'h003EFFD4;
14'd10797:data <=32'h0037FFC3;14'd10798:data <=32'h002CFFB4;14'd10799:data <=32'h001DFFAA;
14'd10800:data <=32'h000CFFA3;14'd10801:data <=32'hFFFAFFA1;14'd10802:data <=32'hFFE9FFA3;
14'd10803:data <=32'hFFD9FFA7;14'd10804:data <=32'hFFCAFFAF;14'd10805:data <=32'hFFBDFFBA;
14'd10806:data <=32'hFFB3FFC8;14'd10807:data <=32'hFFADFFD8;14'd10808:data <=32'hFFABFFE7;
14'd10809:data <=32'hFFADFFF6;14'd10810:data <=32'hFFB30001;14'd10811:data <=32'hFFBA0009;
14'd10812:data <=32'hFFC1000D;14'd10813:data <=32'hFFC6000F;14'd10814:data <=32'hFFC80010;
14'd10815:data <=32'hFFC70011;14'd10816:data <=32'hFFE80004;14'd10817:data <=32'hFFDE0001;
14'd10818:data <=32'hFFD50009;14'd10819:data <=32'hFFC40031;14'd10820:data <=32'hFFB10038;
14'd10821:data <=32'hFFBD0044;14'd10822:data <=32'hFFCA004C;14'd10823:data <=32'hFFD90051;
14'd10824:data <=32'hFFE70052;14'd10825:data <=32'hFFF40052;14'd10826:data <=32'h0001004F;
14'd10827:data <=32'h000C004A;14'd10828:data <=32'h00160042;14'd10829:data <=32'h001E0039;
14'd10830:data <=32'h0023002E;14'd10831:data <=32'h00240023;14'd10832:data <=32'h00210019;
14'd10833:data <=32'h001B0012;14'd10834:data <=32'h00140010;14'd10835:data <=32'h000E0012;
14'd10836:data <=32'h000A0016;14'd10837:data <=32'h000B001C;14'd10838:data <=32'h00100020;
14'd10839:data <=32'h00160023;14'd10840:data <=32'h001E0022;14'd10841:data <=32'h0025001E;
14'd10842:data <=32'h002A0018;14'd10843:data <=32'h002D0011;14'd10844:data <=32'h002F0009;
14'd10845:data <=32'h002E0002;14'd10846:data <=32'h002DFFFB;14'd10847:data <=32'h0029FFF4;
14'd10848:data <=32'h0024FFEF;14'd10849:data <=32'h001DFFEA;14'd10850:data <=32'h0015FFE9;
14'd10851:data <=32'h000DFFEA;14'd10852:data <=32'h0005FFEF;14'd10853:data <=32'h0001FFF7;
14'd10854:data <=32'h00000000;14'd10855:data <=32'h00030008;14'd10856:data <=32'h000A000F;
14'd10857:data <=32'h00140013;14'd10858:data <=32'h001F0012;14'd10859:data <=32'h0029000D;
14'd10860:data <=32'h00310005;14'd10861:data <=32'h0036FFFC;14'd10862:data <=32'h0037FFF2;
14'd10863:data <=32'h0037FFE8;14'd10864:data <=32'h0036FFDE;14'd10865:data <=32'h0033FFD6;
14'd10866:data <=32'h002FFFCE;14'd10867:data <=32'h002AFFC6;14'd10868:data <=32'h0023FFBE;
14'd10869:data <=32'h001BFFB7;14'd10870:data <=32'h0011FFB1;14'd10871:data <=32'h0006FFAD;
14'd10872:data <=32'hFFFAFFAB;14'd10873:data <=32'hFFEFFFAB;14'd10874:data <=32'hFFE5FFAC;
14'd10875:data <=32'hFFDAFFAE;14'd10876:data <=32'hFFCFFFB0;14'd10877:data <=32'hFFC3FFB3;
14'd10878:data <=32'hFFB5FFB8;14'd10879:data <=32'hFFA6FFC1;14'd10880:data <=32'hFFDF0002;
14'd10881:data <=32'hFFDDFFFB;14'd10882:data <=32'hFFD3FFF2;14'd10883:data <=32'hFF92FFE2;
14'd10884:data <=32'hFF75FFF7;14'd10885:data <=32'hFF790012;14'd10886:data <=32'hFF83002B;
14'd10887:data <=32'hFF930040;14'd10888:data <=32'hFFA6004F;14'd10889:data <=32'hFFBA005A;
14'd10890:data <=32'hFFCF005F;14'd10891:data <=32'hFFE40060;14'd10892:data <=32'hFFF8005B;
14'd10893:data <=32'h000A0052;14'd10894:data <=32'h00170045;14'd10895:data <=32'h001F0036;
14'd10896:data <=32'h00220026;14'd10897:data <=32'h001E0017;14'd10898:data <=32'h0016000D;
14'd10899:data <=32'h000D0008;14'd10900:data <=32'h00030008;14'd10901:data <=32'hFFFC000C;
14'd10902:data <=32'hFFF90011;14'd10903:data <=32'hFFF90017;14'd10904:data <=32'hFFFA001D;
14'd10905:data <=32'hFFFF0020;14'd10906:data <=32'h00030022;14'd10907:data <=32'h00070023;
14'd10908:data <=32'h000B0023;14'd10909:data <=32'h00100022;14'd10910:data <=32'h00140021;
14'd10911:data <=32'h0018001E;14'd10912:data <=32'h001C001B;14'd10913:data <=32'h001E0017;
14'd10914:data <=32'h001F0012;14'd10915:data <=32'h001F000D;14'd10916:data <=32'h001D000A;
14'd10917:data <=32'h001A0008;14'd10918:data <=32'h00190008;14'd10919:data <=32'h0019000A;
14'd10920:data <=32'h001A000A;14'd10921:data <=32'h001C000A;14'd10922:data <=32'h001F0008;
14'd10923:data <=32'h00210005;14'd10924:data <=32'h00220001;14'd10925:data <=32'h0021FFFE;
14'd10926:data <=32'h001FFFFB;14'd10927:data <=32'h001CFFFB;14'd10928:data <=32'h001BFFFD;
14'd10929:data <=32'h001B0000;14'd10930:data <=32'h001F0002;14'd10931:data <=32'h00240004;
14'd10932:data <=32'h002C0002;14'd10933:data <=32'h0034FFFD;14'd10934:data <=32'h003BFFF6;
14'd10935:data <=32'h0041FFEC;14'd10936:data <=32'h0044FFDF;14'd10937:data <=32'h0045FFD2;
14'd10938:data <=32'h0044FFC2;14'd10939:data <=32'h003FFFB2;14'd10940:data <=32'h0035FFA1;
14'd10941:data <=32'h0027FF90;14'd10942:data <=32'h0012FF82;14'd10943:data <=32'hFFF8FF79;
14'd10944:data <=32'hFFEAFFC6;14'd10945:data <=32'hFFE1FFBF;14'd10946:data <=32'hFFDEFFB5;
14'd10947:data <=32'hFFD8FF8C;14'd10948:data <=32'hFFA8FF95;14'd10949:data <=32'hFF97FFAA;
14'd10950:data <=32'hFF8DFFC1;14'd10951:data <=32'hFF89FFD9;14'd10952:data <=32'hFF89FFEF;
14'd10953:data <=32'hFF8E0004;14'd10954:data <=32'hFF950016;14'd10955:data <=32'hFFA00026;
14'd10956:data <=32'hFFAE0033;14'd10957:data <=32'hFFBD003C;14'd10958:data <=32'hFFCD003F;
14'd10959:data <=32'hFFDD003F;14'd10960:data <=32'hFFE9003A;14'd10961:data <=32'hFFF20034;
14'd10962:data <=32'hFFF8002E;14'd10963:data <=32'hFFFA0028;14'd10964:data <=32'hFFFB0025;
14'd10965:data <=32'hFFFC0023;14'd10966:data <=32'hFFFE0022;14'd10967:data <=32'h00010021;
14'd10968:data <=32'h0005001E;14'd10969:data <=32'h0007001A;14'd10970:data <=32'h00080015;
14'd10971:data <=32'h00070010;14'd10972:data <=32'h0004000C;14'd10973:data <=32'hFFFF000A;
14'd10974:data <=32'hFFFB000B;14'd10975:data <=32'hFFF7000E;14'd10976:data <=32'hFFF50011;
14'd10977:data <=32'hFFF40016;14'd10978:data <=32'hFFF4001A;14'd10979:data <=32'hFFF6001F;
14'd10980:data <=32'hFFF80024;14'd10981:data <=32'hFFFC0029;14'd10982:data <=32'h0002002D;
14'd10983:data <=32'h00090030;14'd10984:data <=32'h00110031;14'd10985:data <=32'h001C0030;
14'd10986:data <=32'h0025002B;14'd10987:data <=32'h002D0023;14'd10988:data <=32'h00310019;
14'd10989:data <=32'h0032000E;14'd10990:data <=32'h002E0005;14'd10991:data <=32'h0028FFFF;
14'd10992:data <=32'h0021FFFC;14'd10993:data <=32'h001AFFFD;14'd10994:data <=32'h00160001;
14'd10995:data <=32'h00150007;14'd10996:data <=32'h0017000D;14'd10997:data <=32'h001D0011;
14'd10998:data <=32'h00250014;14'd10999:data <=32'h002E0013;14'd11000:data <=32'h00370010;
14'd11001:data <=32'h0041000A;14'd11002:data <=32'h004A0001;14'd11003:data <=32'h0052FFF4;
14'd11004:data <=32'h0058FFE4;14'd11005:data <=32'h0059FFD1;14'd11006:data <=32'h0055FFBC;
14'd11007:data <=32'h004AFFA8;14'd11008:data <=32'h0047FFBF;14'd11009:data <=32'h0041FFA6;
14'd11010:data <=32'h0037FF99;14'd11011:data <=32'h002DFFAA;14'd11012:data <=32'h0004FFA2;
14'd11013:data <=32'hFFF6FFA6;14'd11014:data <=32'hFFEBFFAB;14'd11015:data <=32'hFFE3FFB2;
14'd11016:data <=32'hFFDCFFB7;14'd11017:data <=32'hFFD5FFBC;14'd11018:data <=32'hFFCEFFC2;
14'd11019:data <=32'hFFC7FFC8;14'd11020:data <=32'hFFC1FFD0;14'd11021:data <=32'hFFBCFFDA;
14'd11022:data <=32'hFFB9FFE3;14'd11023:data <=32'hFFB8FFEC;14'd11024:data <=32'hFFB7FFF5;
14'd11025:data <=32'hFFB7FFFD;14'd11026:data <=32'hFFB70006;14'd11027:data <=32'hFFB70010;
14'd11028:data <=32'hFFBA001B;14'd11029:data <=32'hFFC00026;14'd11030:data <=32'hFFCA0031;
14'd11031:data <=32'hFFD70039;14'd11032:data <=32'hFFE6003D;14'd11033:data <=32'hFFF5003B;
14'd11034:data <=32'h00030035;14'd11035:data <=32'h000D002A;14'd11036:data <=32'h0013001E;
14'd11037:data <=32'h00130012;14'd11038:data <=32'h00100008;14'd11039:data <=32'h000AFFFF;
14'd11040:data <=32'h0003FFFA;14'd11041:data <=32'hFFFAFFF7;14'd11042:data <=32'hFFF1FFF7;
14'd11043:data <=32'hFFE9FFFA;14'd11044:data <=32'hFFE10000;14'd11045:data <=32'hFFDB0008;
14'd11046:data <=32'hFFD70012;14'd11047:data <=32'hFFD7001D;14'd11048:data <=32'hFFDA0029;
14'd11049:data <=32'hFFE20033;14'd11050:data <=32'hFFEC003B;14'd11051:data <=32'hFFF8003F;
14'd11052:data <=32'h0003003E;14'd11053:data <=32'h000D003B;14'd11054:data <=32'h00150036;
14'd11055:data <=32'h00190031;14'd11056:data <=32'h001C002C;14'd11057:data <=32'h001D0029;
14'd11058:data <=32'h001F0028;14'd11059:data <=32'h00220028;14'd11060:data <=32'h00270028;
14'd11061:data <=32'h002C0026;14'd11062:data <=32'h00330023;14'd11063:data <=32'h0039001E;
14'd11064:data <=32'h003F0018;14'd11065:data <=32'h00430011;14'd11066:data <=32'h00470009;
14'd11067:data <=32'h004A0001;14'd11068:data <=32'h004CFFF7;14'd11069:data <=32'h004DFFEC;
14'd11070:data <=32'h004CFFE0;14'd11071:data <=32'h0047FFD4;14'd11072:data <=32'h00660017;
14'd11073:data <=32'h0077FFFC;14'd11074:data <=32'h0076FFE0;14'd11075:data <=32'h0031FFD0;
14'd11076:data <=32'h000FFFCA;14'd11077:data <=32'h000AFFD1;14'd11078:data <=32'h0009FFD8;
14'd11079:data <=32'h000BFFDE;14'd11080:data <=32'h000FFFDF;14'd11081:data <=32'h0013FFDC;
14'd11082:data <=32'h0015FFD6;14'd11083:data <=32'h0015FFCF;14'd11084:data <=32'h0011FFC8;
14'd11085:data <=32'h000BFFC0;14'd11086:data <=32'h0002FFBB;14'd11087:data <=32'hFFF8FFB7;
14'd11088:data <=32'hFFECFFB5;14'd11089:data <=32'hFFDFFFB5;14'd11090:data <=32'hFFD0FFB8;
14'd11091:data <=32'hFFC2FFC0;14'd11092:data <=32'hFFB5FFCD;14'd11093:data <=32'hFFABFFDD;
14'd11094:data <=32'hFFA7FFF0;14'd11095:data <=32'hFFA90005;14'd11096:data <=32'hFFB10016;
14'd11097:data <=32'hFFBD0024;14'd11098:data <=32'hFFCD002C;14'd11099:data <=32'hFFDC0030;
14'd11100:data <=32'hFFEA002E;14'd11101:data <=32'hFFF60029;14'd11102:data <=32'hFFFF0022;
14'd11103:data <=32'h0005001A;14'd11104:data <=32'h00070012;14'd11105:data <=32'h0009000A;
14'd11106:data <=32'h00070001;14'd11107:data <=32'h0004FFFA;14'd11108:data <=32'hFFFEFFF4;
14'd11109:data <=32'hFFF7FFF0;14'd11110:data <=32'hFFEDFFEE;14'd11111:data <=32'hFFE4FFF0;
14'd11112:data <=32'hFFDCFFF4;14'd11113:data <=32'hFFD5FFFB;14'd11114:data <=32'hFFD10003;
14'd11115:data <=32'hFFCF000B;14'd11116:data <=32'hFFCE0014;14'd11117:data <=32'hFFCE001B;
14'd11118:data <=32'hFFCF0023;14'd11119:data <=32'hFFD0002B;14'd11120:data <=32'hFFD10035;
14'd11121:data <=32'hFFD50040;14'd11122:data <=32'hFFDC004C;14'd11123:data <=32'hFFE70058;
14'd11124:data <=32'hFFF60061;14'd11125:data <=32'h00090067;14'd11126:data <=32'h001D0068;
14'd11127:data <=32'h00310062;14'd11128:data <=32'h00430059;14'd11129:data <=32'h0053004B;
14'd11130:data <=32'h005E003B;14'd11131:data <=32'h00660029;14'd11132:data <=32'h006A0017;
14'd11133:data <=32'h006A0004;14'd11134:data <=32'h0067FFF0;14'd11135:data <=32'h005EFFDF;
14'd11136:data <=32'h0036003A;14'd11137:data <=32'h004D0032;14'd11138:data <=32'h0060001C;
14'd11139:data <=32'h0050FFD5;14'd11140:data <=32'h0027FFCA;14'd11141:data <=32'h001AFFCF;
14'd11142:data <=32'h0012FFD8;14'd11143:data <=32'h000FFFE1;14'd11144:data <=32'h0011FFE8;
14'd11145:data <=32'h0015FFEC;14'd11146:data <=32'h001AFFED;14'd11147:data <=32'h001EFFEA;
14'd11148:data <=32'h0021FFE5;14'd11149:data <=32'h0022FFDF;14'd11150:data <=32'h0021FFD9;
14'd11151:data <=32'h001FFFD2;14'd11152:data <=32'h001BFFCA;14'd11153:data <=32'h0014FFC3;
14'd11154:data <=32'h000BFFBD;14'd11155:data <=32'hFFFFFFB9;14'd11156:data <=32'hFFF2FFB9;
14'd11157:data <=32'hFFE4FFBC;14'd11158:data <=32'hFFD9FFC4;14'd11159:data <=32'hFFD0FFCF;
14'd11160:data <=32'hFFCCFFDC;14'd11161:data <=32'hFFCBFFE7;14'd11162:data <=32'hFFCEFFF1;
14'd11163:data <=32'hFFD1FFF8;14'd11164:data <=32'hFFD6FFFD;14'd11165:data <=32'hFFDA0001;
14'd11166:data <=32'hFFDD0004;14'd11167:data <=32'hFFE00006;14'd11168:data <=32'hFFE40009;
14'd11169:data <=32'hFFE8000B;14'd11170:data <=32'hFFED000D;14'd11171:data <=32'hFFF2000C;
14'd11172:data <=32'hFFF8000A;14'd11173:data <=32'hFFFC0006;14'd11174:data <=32'hFFFE0001;
14'd11175:data <=32'hFFFFFFFB;14'd11176:data <=32'hFFFDFFF5;14'd11177:data <=32'hFFFAFFEF;
14'd11178:data <=32'hFFF5FFEB;14'd11179:data <=32'hFFEFFFE6;14'd11180:data <=32'hFFE8FFE3;
14'd11181:data <=32'hFFDEFFE1;14'd11182:data <=32'hFFD2FFE1;14'd11183:data <=32'hFFC5FFE5;
14'd11184:data <=32'hFFB7FFEE;14'd11185:data <=32'hFFAAFFFB;14'd11186:data <=32'hFFA1000E;
14'd11187:data <=32'hFF9D0024;14'd11188:data <=32'hFFA0003D;14'd11189:data <=32'hFFAB0055;
14'd11190:data <=32'hFFBC0068;14'd11191:data <=32'hFFD10077;14'd11192:data <=32'hFFEA0080;
14'd11193:data <=32'h00030082;14'd11194:data <=32'h001C007F;14'd11195:data <=32'h00320077;
14'd11196:data <=32'h0047006A;14'd11197:data <=32'h00570059;14'd11198:data <=32'h00640045;
14'd11199:data <=32'h006B0030;14'd11200:data <=32'h00320038;14'd11201:data <=32'h00400035;
14'd11202:data <=32'h00520031;14'd11203:data <=32'h006C0025;14'd11204:data <=32'h0050000D;
14'd11205:data <=32'h004A0005;14'd11206:data <=32'h00460000;14'd11207:data <=32'h0043FFFC;
14'd11208:data <=32'h0043FFF8;14'd11209:data <=32'h0042FFF2;14'd11210:data <=32'h0041FFEB;
14'd11211:data <=32'h003FFFE3;14'd11212:data <=32'h003AFFDA;14'd11213:data <=32'h0033FFD4;
14'd11214:data <=32'h002AFFCF;14'd11215:data <=32'h0022FFCC;14'd11216:data <=32'h001BFFCB;
14'd11217:data <=32'h0013FFCB;14'd11218:data <=32'h000DFFCB;14'd11219:data <=32'h0006FFCD;
14'd11220:data <=32'hFFFEFFCF;14'd11221:data <=32'hFFF8FFD3;14'd11222:data <=32'hFFF4FFD9;
14'd11223:data <=32'hFFF1FFE0;14'd11224:data <=32'hFFF2FFE7;14'd11225:data <=32'hFFF5FFEC;
14'd11226:data <=32'hFFF9FFEF;14'd11227:data <=32'hFFFEFFEE;14'd11228:data <=32'h0001FFEA;
14'd11229:data <=32'h0001FFE6;14'd11230:data <=32'hFFFEFFE1;14'd11231:data <=32'hFFF8FFDE;
14'd11232:data <=32'hFFF2FFDE;14'd11233:data <=32'hFFECFFE0;14'd11234:data <=32'hFFE7FFE5;
14'd11235:data <=32'hFFE5FFEA;14'd11236:data <=32'hFFE5FFF0;14'd11237:data <=32'hFFE7FFF5;
14'd11238:data <=32'hFFE9FFF8;14'd11239:data <=32'hFFEDFFFA;14'd11240:data <=32'hFFF1FFFB;
14'd11241:data <=32'hFFF5FFFA;14'd11242:data <=32'hFFF8FFF8;14'd11243:data <=32'hFFFBFFF3;
14'd11244:data <=32'hFFFCFFED;14'd11245:data <=32'hFFFBFFE6;14'd11246:data <=32'hFFF6FFDD;
14'd11247:data <=32'hFFEDFFD6;14'd11248:data <=32'hFFE1FFD1;14'd11249:data <=32'hFFD2FFD0;
14'd11250:data <=32'hFFC1FFD5;14'd11251:data <=32'hFFB2FFE0;14'd11252:data <=32'hFFA6FFF0;
14'd11253:data <=32'hFFA00002;14'd11254:data <=32'hFF9F0015;14'd11255:data <=32'hFFA20028;
14'd11256:data <=32'hFFAA0039;14'd11257:data <=32'hFFB50047;14'd11258:data <=32'hFFC10052;
14'd11259:data <=32'hFFCF005B;14'd11260:data <=32'hFFDD0061;14'd11261:data <=32'hFFEC0065;
14'd11262:data <=32'hFFFC0066;14'd11263:data <=32'h000C0064;14'd11264:data <=32'h001C006A;
14'd11265:data <=32'h00300067;14'd11266:data <=32'h00390062;14'd11267:data <=32'h00160068;
14'd11268:data <=32'h000A005C;14'd11269:data <=32'h0016005E;14'd11270:data <=32'h0024005F;
14'd11271:data <=32'h0033005D;14'd11272:data <=32'h00450057;14'd11273:data <=32'h0056004B;
14'd11274:data <=32'h0065003B;14'd11275:data <=32'h006F0026;14'd11276:data <=32'h0073000F;
14'd11277:data <=32'h0070FFF8;14'd11278:data <=32'h0068FFE3;14'd11279:data <=32'h005CFFD2;
14'd11280:data <=32'h004DFFC6;14'd11281:data <=32'h003CFFBE;14'd11282:data <=32'h002BFFB9;
14'd11283:data <=32'h001BFFB9;14'd11284:data <=32'h000AFFBC;14'd11285:data <=32'hFFFCFFC3;
14'd11286:data <=32'hFFF1FFCE;14'd11287:data <=32'hFFEAFFDB;14'd11288:data <=32'hFFE8FFE9;
14'd11289:data <=32'hFFEBFFF6;14'd11290:data <=32'hFFF20000;14'd11291:data <=32'hFFFD0006;
14'd11292:data <=32'h00080007;14'd11293:data <=32'h00110003;14'd11294:data <=32'h0017FFFC;
14'd11295:data <=32'h001AFFF4;14'd11296:data <=32'h0019FFED;14'd11297:data <=32'h0017FFE7;
14'd11298:data <=32'h0013FFE2;14'd11299:data <=32'h000FFFE0;14'd11300:data <=32'h000BFFDE;
14'd11301:data <=32'h0009FFDC;14'd11302:data <=32'h0005FFDB;14'd11303:data <=32'h0001FFDA;
14'd11304:data <=32'hFFFEFFDA;14'd11305:data <=32'hFFFAFFDA;14'd11306:data <=32'hFFF7FFDB;
14'd11307:data <=32'hFFF5FFDB;14'd11308:data <=32'hFFF2FFDC;14'd11309:data <=32'hFFF0FFDB;
14'd11310:data <=32'hFFEEFFDA;14'd11311:data <=32'hFFEBFFD8;14'd11312:data <=32'hFFE5FFD6;
14'd11313:data <=32'hFFDEFFD6;14'd11314:data <=32'hFFD5FFD8;14'd11315:data <=32'hFFCDFFDE;
14'd11316:data <=32'hFFC7FFE5;14'd11317:data <=32'hFFC3FFEF;14'd11318:data <=32'hFFC2FFF7;
14'd11319:data <=32'hFFC4FFFF;14'd11320:data <=32'hFFC70005;14'd11321:data <=32'hFFCA0009;
14'd11322:data <=32'hFFCB000B;14'd11323:data <=32'hFFCB000D;14'd11324:data <=32'hFFC90010;
14'd11325:data <=32'hFFC60014;14'd11326:data <=32'hFFC4001A;14'd11327:data <=32'hFFC30022;
14'd11328:data <=32'hFFC1005F;14'd11329:data <=32'hFFD1006C;14'd11330:data <=32'hFFE00069;
14'd11331:data <=32'hFFC80034;14'd11332:data <=32'hFFB10035;14'd11333:data <=32'hFFB40047;
14'd11334:data <=32'hFFBE005B;14'd11335:data <=32'hFFCC006C;14'd11336:data <=32'hFFE2007A;
14'd11337:data <=32'hFFFB0082;14'd11338:data <=32'h00180082;14'd11339:data <=32'h0033007A;
14'd11340:data <=32'h004A006B;14'd11341:data <=32'h005C0057;14'd11342:data <=32'h00670041;
14'd11343:data <=32'h006C002A;14'd11344:data <=32'h006C0013;14'd11345:data <=32'h0067FFFF;
14'd11346:data <=32'h005FFFED;14'd11347:data <=32'h0053FFDE;14'd11348:data <=32'h0045FFD3;
14'd11349:data <=32'h0035FFCB;14'd11350:data <=32'h0024FFC8;14'd11351:data <=32'h0014FFCA;
14'd11352:data <=32'h0006FFD2;14'd11353:data <=32'hFFFDFFDB;14'd11354:data <=32'hFFF8FFE6;
14'd11355:data <=32'hFFF7FFF0;14'd11356:data <=32'hFFFAFFF9;14'd11357:data <=32'hFFFDFFFF;
14'd11358:data <=32'h00020002;14'd11359:data <=32'h00060004;14'd11360:data <=32'h00090005;
14'd11361:data <=32'h000D0006;14'd11362:data <=32'h00110007;14'd11363:data <=32'h00160008;
14'd11364:data <=32'h001C0007;14'd11365:data <=32'h00230004;14'd11366:data <=32'h002AFFFE;
14'd11367:data <=32'h002FFFF6;14'd11368:data <=32'h0031FFEC;14'd11369:data <=32'h0031FFE1;
14'd11370:data <=32'h002EFFD6;14'd11371:data <=32'h0029FFCC;14'd11372:data <=32'h0022FFC3;
14'd11373:data <=32'h0018FFBC;14'd11374:data <=32'h000EFFB6;14'd11375:data <=32'h0001FFB2;
14'd11376:data <=32'hFFF4FFB0;14'd11377:data <=32'hFFE6FFB2;14'd11378:data <=32'hFFD7FFB8;
14'd11379:data <=32'hFFCBFFC2;14'd11380:data <=32'hFFC2FFCE;14'd11381:data <=32'hFFBDFFDD;
14'd11382:data <=32'hFFBEFFEC;14'd11383:data <=32'hFFC3FFF8;14'd11384:data <=32'hFFCB0001;
14'd11385:data <=32'hFFD40005;14'd11386:data <=32'hFFDD0004;14'd11387:data <=32'hFFE20000;
14'd11388:data <=32'hFFE4FFFB;14'd11389:data <=32'hFFE1FFF5;14'd11390:data <=32'hFFDDFFF2;
14'd11391:data <=32'hFFD6FFF0;14'd11392:data <=32'hFFB30000;14'd11393:data <=32'hFFAD000C;
14'd11394:data <=32'hFFB30016;14'd11395:data <=32'hFFD20005;14'd11396:data <=32'hFFB5FFFD;
14'd11397:data <=32'hFFAD000A;14'd11398:data <=32'hFFAA001A;14'd11399:data <=32'hFFAA002B;
14'd11400:data <=32'hFFB0003E;14'd11401:data <=32'hFFBD004E;14'd11402:data <=32'hFFCD005A;
14'd11403:data <=32'hFFE00061;14'd11404:data <=32'hFFF30062;14'd11405:data <=32'h0004005F;
14'd11406:data <=32'h00120059;14'd11407:data <=32'h001E0051;14'd11408:data <=32'h00270048;
14'd11409:data <=32'h002E003F;14'd11410:data <=32'h00340036;14'd11411:data <=32'h0038002C;
14'd11412:data <=32'h003B0021;14'd11413:data <=32'h003C0017;14'd11414:data <=32'h003A000D;
14'd11415:data <=32'h00360004;14'd11416:data <=32'h0031FFFD;14'd11417:data <=32'h002BFFF9;
14'd11418:data <=32'h0026FFF6;14'd11419:data <=32'h0022FFF3;14'd11420:data <=32'h001EFFF1;
14'd11421:data <=32'h0019FFEE;14'd11422:data <=32'h0014FFED;14'd11423:data <=32'h000DFFEC;
14'd11424:data <=32'h0006FFEE;14'd11425:data <=32'hFFFFFFF3;14'd11426:data <=32'hFFF9FFFB;
14'd11427:data <=32'hFFF80005;14'd11428:data <=32'hFFFA0010;14'd11429:data <=32'h0001001A;
14'd11430:data <=32'h000B0021;14'd11431:data <=32'h00180024;14'd11432:data <=32'h00260022;
14'd11433:data <=32'h0033001C;14'd11434:data <=32'h003E0013;14'd11435:data <=32'h00470006;
14'd11436:data <=32'h004CFFF8;14'd11437:data <=32'h004DFFE9;14'd11438:data <=32'h004CFFD8;
14'd11439:data <=32'h0047FFC8;14'd11440:data <=32'h003DFFB9;14'd11441:data <=32'h002FFFAD;
14'd11442:data <=32'h001EFFA4;14'd11443:data <=32'h000CFFA1;14'd11444:data <=32'hFFF9FFA3;
14'd11445:data <=32'hFFE9FFAA;14'd11446:data <=32'hFFDDFFB4;14'd11447:data <=32'hFFD5FFC0;
14'd11448:data <=32'hFFD2FFCC;14'd11449:data <=32'hFFD2FFD5;14'd11450:data <=32'hFFD4FFDB;
14'd11451:data <=32'hFFD6FFDE;14'd11452:data <=32'hFFD6FFE0;14'd11453:data <=32'hFFD5FFE1;
14'd11454:data <=32'hFFD3FFE2;14'd11455:data <=32'hFFCFFFE4;14'd11456:data <=32'hFFEFFFE7;
14'd11457:data <=32'hFFE7FFDE;14'd11458:data <=32'hFFDDFFDF;14'd11459:data <=32'hFFC4FFFB;
14'd11460:data <=32'hFFACFFF6;14'd11461:data <=32'hFFAB0002;14'd11462:data <=32'hFFAD000E;
14'd11463:data <=32'hFFB0001B;14'd11464:data <=32'hFFB70027;14'd11465:data <=32'hFFC10032;
14'd11466:data <=32'hFFCE0038;14'd11467:data <=32'hFFDB003B;14'd11468:data <=32'hFFE80039;
14'd11469:data <=32'hFFF10034;14'd11470:data <=32'hFFF7002D;14'd11471:data <=32'hFFF90028;
14'd11472:data <=32'hFFF80023;14'd11473:data <=32'hFFF60022;14'd11474:data <=32'hFFF50024;
14'd11475:data <=32'hFFF50026;14'd11476:data <=32'hFFF70029;14'd11477:data <=32'hFFFB002C;
14'd11478:data <=32'hFFFF002F;14'd11479:data <=32'h00040030;14'd11480:data <=32'h000A0030;
14'd11481:data <=32'h00110030;14'd11482:data <=32'h0018002E;14'd11483:data <=32'h0020002B;
14'd11484:data <=32'h00270024;14'd11485:data <=32'h002C001B;14'd11486:data <=32'h002E0010;
14'd11487:data <=32'h002D0005;14'd11488:data <=32'h0027FFFB;14'd11489:data <=32'h001EFFF4;
14'd11490:data <=32'h0013FFF1;14'd11491:data <=32'h0008FFF3;14'd11492:data <=32'hFFFFFFF9;
14'd11493:data <=32'hFFFA0001;14'd11494:data <=32'hFFF9000C;14'd11495:data <=32'hFFFB0015;
14'd11496:data <=32'h0001001D;14'd11497:data <=32'h00090022;14'd11498:data <=32'h00120026;
14'd11499:data <=32'h001C0027;14'd11500:data <=32'h00250026;14'd11501:data <=32'h00300022;
14'd11502:data <=32'h0039001C;14'd11503:data <=32'h00420014;14'd11504:data <=32'h00480008;
14'd11505:data <=32'h004CFFFC;14'd11506:data <=32'h004DFFEF;14'd11507:data <=32'h004AFFE2;
14'd11508:data <=32'h0045FFD6;14'd11509:data <=32'h003EFFCD;14'd11510:data <=32'h0037FFC6;
14'd11511:data <=32'h0030FFC1;14'd11512:data <=32'h002BFFBC;14'd11513:data <=32'h0025FFB5;
14'd11514:data <=32'h001EFFAE;14'd11515:data <=32'h0015FFA7;14'd11516:data <=32'h0009FF9F;
14'd11517:data <=32'hFFFAFF9A;14'd11518:data <=32'hFFE8FF99;14'd11519:data <=32'hFFD6FF9C;
14'd11520:data <=32'hFFF6FFF2;14'd11521:data <=32'hFFFAFFE8;14'd11522:data <=32'hFFF7FFD8;
14'd11523:data <=32'hFFBDFFB2;14'd11524:data <=32'hFF9BFFB4;14'd11525:data <=32'hFF91FFC9;
14'd11526:data <=32'hFF8CFFE0;14'd11527:data <=32'hFF8CFFF7;14'd11528:data <=32'hFF92000E;
14'd11529:data <=32'hFF9E0022;14'd11530:data <=32'hFFAF0031;14'd11531:data <=32'hFFC2003A;
14'd11532:data <=32'hFFD6003C;14'd11533:data <=32'hFFE70038;14'd11534:data <=32'hFFF4002E;
14'd11535:data <=32'hFFFC0024;14'd11536:data <=32'hFFFD0019;14'd11537:data <=32'hFFFB0010;
14'd11538:data <=32'hFFF7000B;14'd11539:data <=32'hFFF10009;14'd11540:data <=32'hFFED0009;
14'd11541:data <=32'hFFE9000C;14'd11542:data <=32'hFFE6000F;14'd11543:data <=32'hFFE40014;
14'd11544:data <=32'hFFE3001A;14'd11545:data <=32'hFFE40020;14'd11546:data <=32'hFFE70027;
14'd11547:data <=32'hFFED002C;14'd11548:data <=32'hFFF50030;14'd11549:data <=32'hFFFE0031;
14'd11550:data <=32'h0007002F;14'd11551:data <=32'h000F002A;14'd11552:data <=32'h00130023;
14'd11553:data <=32'h0015001C;14'd11554:data <=32'h00130016;14'd11555:data <=32'h00110012;
14'd11556:data <=32'h000E0011;14'd11557:data <=32'h000B0011;14'd11558:data <=32'h000A0012;
14'd11559:data <=32'h000A0014;14'd11560:data <=32'h000B0014;14'd11561:data <=32'h000D0014;
14'd11562:data <=32'h000E0014;14'd11563:data <=32'h000D0013;14'd11564:data <=32'h000D0014;
14'd11565:data <=32'h000D0016;14'd11566:data <=32'h000D0018;14'd11567:data <=32'h000F001C;
14'd11568:data <=32'h0013001F;14'd11569:data <=32'h00180022;14'd11570:data <=32'h001E0023;
14'd11571:data <=32'h00250024;14'd11572:data <=32'h002D0023;14'd11573:data <=32'h00350022;
14'd11574:data <=32'h003F001F;14'd11575:data <=32'h004A001A;14'd11576:data <=32'h00560012;
14'd11577:data <=32'h00620004;14'd11578:data <=32'h006BFFF2;14'd11579:data <=32'h0070FFDB;
14'd11580:data <=32'h006EFFC2;14'd11581:data <=32'h0065FFA9;14'd11582:data <=32'h0054FF92;
14'd11583:data <=32'h003DFF81;14'd11584:data <=32'h000DFFCE;14'd11585:data <=32'h000EFFC6;
14'd11586:data <=32'h0015FFBA;14'd11587:data <=32'h001EFF88;14'd11588:data <=32'hFFF1FF78;
14'd11589:data <=32'hFFD9FF80;14'd11590:data <=32'hFFC3FF8D;14'd11591:data <=32'hFFB1FF9E;
14'd11592:data <=32'hFFA4FFB3;14'd11593:data <=32'hFF9DFFCA;14'd11594:data <=32'hFF9DFFE1;
14'd11595:data <=32'hFFA3FFF5;14'd11596:data <=32'hFFAD0004;14'd11597:data <=32'hFFB9000F;
14'd11598:data <=32'hFFC50014;14'd11599:data <=32'hFFCF0015;14'd11600:data <=32'hFFD60015;
14'd11601:data <=32'hFFDB0014;14'd11602:data <=32'hFFDE0013;14'd11603:data <=32'hFFE10014;
14'd11604:data <=32'hFFE40015;14'd11605:data <=32'hFFE80014;14'd11606:data <=32'hFFEB0014;
14'd11607:data <=32'hFFED0012;14'd11608:data <=32'hFFEF0010;14'd11609:data <=32'hFFEF000F;
14'd11610:data <=32'hFFEF000E;14'd11611:data <=32'hFFEE000E;14'd11612:data <=32'hFFEE000F;
14'd11613:data <=32'hFFEE0010;14'd11614:data <=32'hFFEF0010;14'd11615:data <=32'hFFEF000F;
14'd11616:data <=32'hFFEE000F;14'd11617:data <=32'hFFEC000F;14'd11618:data <=32'hFFEA0011;
14'd11619:data <=32'hFFE70015;14'd11620:data <=32'hFFE6001B;14'd11621:data <=32'hFFE80022;
14'd11622:data <=32'hFFEC0029;14'd11623:data <=32'hFFF3002E;14'd11624:data <=32'hFFFC0031;
14'd11625:data <=32'h00050030;14'd11626:data <=32'h000C002C;14'd11627:data <=32'h00120026;
14'd11628:data <=32'h0014001F;14'd11629:data <=32'h00140019;14'd11630:data <=32'h00110015;
14'd11631:data <=32'h000E0012;14'd11632:data <=32'h000A0012;14'd11633:data <=32'h00060014;
14'd11634:data <=32'h00030018;14'd11635:data <=32'h0002001D;14'd11636:data <=32'h00030024;
14'd11637:data <=32'h0005002C;14'd11638:data <=32'h000C0034;14'd11639:data <=32'h0016003D;
14'd11640:data <=32'h00240042;14'd11641:data <=32'h00360043;14'd11642:data <=32'h004A003E;
14'd11643:data <=32'h005E0033;14'd11644:data <=32'h006E0020;14'd11645:data <=32'h0078000A;
14'd11646:data <=32'h007CFFF0;14'd11647:data <=32'h0078FFD7;14'd11648:data <=32'h005CFFEB;
14'd11649:data <=32'h0063FFD7;14'd11650:data <=32'h0065FFCC;14'd11651:data <=32'h0062FFD3;
14'd11652:data <=32'h0044FFB6;14'd11653:data <=32'h0037FFAE;14'd11654:data <=32'h002AFFA8;
14'd11655:data <=32'h001CFFA5;14'd11656:data <=32'h000EFFA4;14'd11657:data <=32'h0000FFA7;
14'd11658:data <=32'hFFF5FFAB;14'd11659:data <=32'hFFECFFB1;14'd11660:data <=32'hFFE5FFB7;
14'd11661:data <=32'hFFE0FFBC;14'd11662:data <=32'hFFDAFFC0;14'd11663:data <=32'hFFD4FFC3;
14'd11664:data <=32'hFFCCFFC9;14'd11665:data <=32'hFFC4FFCF;14'd11666:data <=32'hFFBCFFDA;
14'd11667:data <=32'hFFB7FFE7;14'd11668:data <=32'hFFB6FFF5;14'd11669:data <=32'hFFB90004;
14'd11670:data <=32'hFFC00010;14'd11671:data <=32'hFFCA001A;14'd11672:data <=32'hFFD5001F;
14'd11673:data <=32'hFFE00022;14'd11674:data <=32'hFFEA0021;14'd11675:data <=32'hFFF3001E;
14'd11676:data <=32'hFFFB0019;14'd11677:data <=32'h00010012;14'd11678:data <=32'h0005000A;
14'd11679:data <=32'h00050002;14'd11680:data <=32'h0003FFF8;14'd11681:data <=32'hFFFCFFF1;
14'd11682:data <=32'hFFF3FFEB;14'd11683:data <=32'hFFE8FFEA;14'd11684:data <=32'hFFDDFFED;
14'd11685:data <=32'hFFD3FFF5;14'd11686:data <=32'hFFCD0000;14'd11687:data <=32'hFFCB000C;
14'd11688:data <=32'hFFCD0017;14'd11689:data <=32'hFFD30021;14'd11690:data <=32'hFFD90028;
14'd11691:data <=32'hFFE1002C;14'd11692:data <=32'hFFE8002D;14'd11693:data <=32'hFFEE002D;
14'd11694:data <=32'hFFF2002D;14'd11695:data <=32'hFFF5002C;14'd11696:data <=32'hFFF8002C;
14'd11697:data <=32'hFFFB002D;14'd11698:data <=32'hFFFD002D;14'd11699:data <=32'h0000002E;
14'd11700:data <=32'h0002002F;14'd11701:data <=32'h00040031;14'd11702:data <=32'h00070034;
14'd11703:data <=32'h000B0039;14'd11704:data <=32'h0013003D;14'd11705:data <=32'h001D0040;
14'd11706:data <=32'h00280040;14'd11707:data <=32'h0036003C;14'd11708:data <=32'h00420035;
14'd11709:data <=32'h004D0029;14'd11710:data <=32'h0053001B;14'd11711:data <=32'h0054000D;
14'd11712:data <=32'h0053004B;14'd11713:data <=32'h006D003E;14'd11714:data <=32'h0079002A;
14'd11715:data <=32'h00460009;14'd11716:data <=32'h0030FFF5;14'd11717:data <=32'h002FFFF5;
14'd11718:data <=32'h0030FFF5;14'd11719:data <=32'h0031FFF3;14'd11720:data <=32'h0033FFF0;
14'd11721:data <=32'h0035FFEC;14'd11722:data <=32'h0037FFE6;14'd11723:data <=32'h0039FFE0;
14'd11724:data <=32'h003AFFD7;14'd11725:data <=32'h0038FFCC;14'd11726:data <=32'h0034FFBF;
14'd11727:data <=32'h002CFFB2;14'd11728:data <=32'h001EFFA6;14'd11729:data <=32'h000CFF9E;
14'd11730:data <=32'hFFF8FF9C;14'd11731:data <=32'hFFE3FFA0;14'd11732:data <=32'hFFD0FFAB;
14'd11733:data <=32'hFFC2FFBA;14'd11734:data <=32'hFFB9FFCB;14'd11735:data <=32'hFFB6FFDD;
14'd11736:data <=32'hFFB7FFEE;14'd11737:data <=32'hFFBCFFFD;14'd11738:data <=32'hFFC4000A;
14'd11739:data <=32'hFFCD0014;14'd11740:data <=32'hFFD9001A;14'd11741:data <=32'hFFE5001D;
14'd11742:data <=32'hFFF1001C;14'd11743:data <=32'hFFFC0018;14'd11744:data <=32'h00060010;
14'd11745:data <=32'h000B0006;14'd11746:data <=32'h000DFFFA;14'd11747:data <=32'h000AFFF0;
14'd11748:data <=32'h0003FFE7;14'd11749:data <=32'hFFFBFFE2;14'd11750:data <=32'hFFF2FFE0;
14'd11751:data <=32'hFFE9FFE1;14'd11752:data <=32'hFFE1FFE3;14'd11753:data <=32'hFFDBFFE7;
14'd11754:data <=32'hFFD6FFEA;14'd11755:data <=32'hFFD1FFEE;14'd11756:data <=32'hFFCCFFF2;
14'd11757:data <=32'hFFC6FFF7;14'd11758:data <=32'hFFC0FFFF;14'd11759:data <=32'hFFBB0009;
14'd11760:data <=32'hFFB70015;14'd11761:data <=32'hFFB70023;14'd11762:data <=32'hFFBB0030;
14'd11763:data <=32'hFFC1003D;14'd11764:data <=32'hFFCA0049;14'd11765:data <=32'hFFD60053;
14'd11766:data <=32'hFFE2005A;14'd11767:data <=32'hFFF10060;14'd11768:data <=32'h00000063;
14'd11769:data <=32'h00110063;14'd11770:data <=32'h0022005F;14'd11771:data <=32'h00330057;
14'd11772:data <=32'h0042004A;14'd11773:data <=32'h004C003A;14'd11774:data <=32'h00510027;
14'd11775:data <=32'h004F0015;14'd11776:data <=32'h000A0058;14'd11777:data <=32'h00200060;
14'd11778:data <=32'h003A0059;14'd11779:data <=32'h00440012;14'd11780:data <=32'h002AFFFC;
14'd11781:data <=32'h0023FFFE;14'd11782:data <=32'h001E0001;14'd11783:data <=32'h001E0006;
14'd11784:data <=32'h001F0009;14'd11785:data <=32'h0022000C;14'd11786:data <=32'h0026000E;
14'd11787:data <=32'h002E000E;14'd11788:data <=32'h0036000C;14'd11789:data <=32'h003F0006;
14'd11790:data <=32'h0046FFFB;14'd11791:data <=32'h004BFFED;14'd11792:data <=32'h004AFFDD;
14'd11793:data <=32'h0044FFCD;14'd11794:data <=32'h0039FFBF;14'd11795:data <=32'h002AFFB5;
14'd11796:data <=32'h001AFFB1;14'd11797:data <=32'h000AFFB1;14'd11798:data <=32'hFFFCFFB5;
14'd11799:data <=32'hFFF1FFBC;14'd11800:data <=32'hFFE8FFC4;14'd11801:data <=32'hFFE2FFCC;
14'd11802:data <=32'hFFDDFFD4;14'd11803:data <=32'hFFDAFFDD;14'd11804:data <=32'hFFD9FFE6;
14'd11805:data <=32'hFFD9FFEE;14'd11806:data <=32'hFFDCFFF7;14'd11807:data <=32'hFFE1FFFE;
14'd11808:data <=32'hFFE70003;14'd11809:data <=32'hFFEE0004;14'd11810:data <=32'hFFF50004;
14'd11811:data <=32'hFFFA0002;14'd11812:data <=32'hFFFEFFFF;14'd11813:data <=32'h0001FFFC;
14'd11814:data <=32'h0004FFF9;14'd11815:data <=32'h0006FFF5;14'd11816:data <=32'h0007FFF0;
14'd11817:data <=32'h0009FFE9;14'd11818:data <=32'h0009FFE1;14'd11819:data <=32'h0005FFD7;
14'd11820:data <=32'hFFFEFFCD;14'd11821:data <=32'hFFF3FFC5;14'd11822:data <=32'hFFE3FFBF;
14'd11823:data <=32'hFFD1FFBE;14'd11824:data <=32'hFFBFFFC3;14'd11825:data <=32'hFFADFFCE;
14'd11826:data <=32'hFF9EFFDE;14'd11827:data <=32'hFF94FFF1;14'd11828:data <=32'hFF8E0007;
14'd11829:data <=32'hFF8E001D;14'd11830:data <=32'hFF930033;14'd11831:data <=32'hFF9C0049;
14'd11832:data <=32'hFFAA005C;14'd11833:data <=32'hFFBD006C;14'd11834:data <=32'hFFD30077;
14'd11835:data <=32'hFFEC007C;14'd11836:data <=32'h0006007A;14'd11837:data <=32'h001D0071;
14'd11838:data <=32'h00300063;14'd11839:data <=32'h003D0051;14'd11840:data <=32'h00000040;
14'd11841:data <=32'h00070047;14'd11842:data <=32'h00160051;14'd11843:data <=32'h00390050;
14'd11844:data <=32'h002B0034;14'd11845:data <=32'h002C002F;14'd11846:data <=32'h002E002B;
14'd11847:data <=32'h00310027;14'd11848:data <=32'h00330021;14'd11849:data <=32'h0035001D;
14'd11850:data <=32'h00360018;14'd11851:data <=32'h00370013;14'd11852:data <=32'h0039000F;
14'd11853:data <=32'h003B000A;14'd11854:data <=32'h003D0003;14'd11855:data <=32'h003EFFFB;
14'd11856:data <=32'h003DFFF2;14'd11857:data <=32'h0039FFE8;14'd11858:data <=32'h0032FFE0;
14'd11859:data <=32'h0029FFDB;14'd11860:data <=32'h0020FFD9;14'd11861:data <=32'h0018FFDB;
14'd11862:data <=32'h0012FFDE;14'd11863:data <=32'h000FFFE2;14'd11864:data <=32'h000EFFE6;
14'd11865:data <=32'h000FFFE7;14'd11866:data <=32'h0010FFE6;14'd11867:data <=32'h000FFFE4;
14'd11868:data <=32'h000EFFE1;14'd11869:data <=32'h000BFFDF;14'd11870:data <=32'h0007FFDE;
14'd11871:data <=32'h0003FFDF;14'd11872:data <=32'hFFFFFFDF;14'd11873:data <=32'hFFFCFFE1;
14'd11874:data <=32'hFFF9FFE3;14'd11875:data <=32'hFFF7FFE5;14'd11876:data <=32'hFFF4FFE9;
14'd11877:data <=32'hFFF3FFED;14'd11878:data <=32'hFFF3FFF2;14'd11879:data <=32'hFFF6FFF8;
14'd11880:data <=32'hFFFBFFFC;14'd11881:data <=32'h0003FFFD;14'd11882:data <=32'h000CFFFB;
14'd11883:data <=32'h0014FFF4;14'd11884:data <=32'h0019FFE9;14'd11885:data <=32'h001AFFDC;
14'd11886:data <=32'h0017FFCE;14'd11887:data <=32'h000DFFC0;14'd11888:data <=32'hFFFFFFB7;
14'd11889:data <=32'hFFEEFFB2;14'd11890:data <=32'hFFDCFFB1;14'd11891:data <=32'hFFCAFFB5;
14'd11892:data <=32'hFFBBFFBD;14'd11893:data <=32'hFFACFFC8;14'd11894:data <=32'hFFA0FFD7;
14'd11895:data <=32'hFF97FFE8;14'd11896:data <=32'hFF93FFFA;14'd11897:data <=32'hFF92000E;
14'd11898:data <=32'hFF950022;14'd11899:data <=32'hFF9E0035;14'd11900:data <=32'hFFAB0044;
14'd11901:data <=32'hFFBA004F;14'd11902:data <=32'hFFCA0055;14'd11903:data <=32'hFFD80056;
14'd11904:data <=32'hFFE70058;14'd11905:data <=32'hFFF2005B;14'd11906:data <=32'hFFF6005D;
14'd11907:data <=32'hFFD50062;14'd11908:data <=32'hFFCE0057;14'd11909:data <=32'hFFDA0061;
14'd11910:data <=32'hFFEA0069;14'd11911:data <=32'hFFFC006E;14'd11912:data <=32'h0010006E;
14'd11913:data <=32'h00230068;14'd11914:data <=32'h0034005F;14'd11915:data <=32'h00430053;
14'd11916:data <=32'h004E0045;14'd11917:data <=32'h00560034;14'd11918:data <=32'h005B0023;
14'd11919:data <=32'h005C0011;14'd11920:data <=32'h0059FFFE;14'd11921:data <=32'h0051FFEE;
14'd11922:data <=32'h0044FFE0;14'd11923:data <=32'h0035FFD7;14'd11924:data <=32'h0024FFD4;
14'd11925:data <=32'h0014FFD6;14'd11926:data <=32'h0008FFDE;14'd11927:data <=32'h0001FFE8;
14'd11928:data <=32'hFFFEFFF3;14'd11929:data <=32'h0000FFFC;14'd11930:data <=32'h00050003;
14'd11931:data <=32'h000B0007;14'd11932:data <=32'h00110007;14'd11933:data <=32'h00170006;
14'd11934:data <=32'h001B0003;14'd11935:data <=32'h001EFFFF;14'd11936:data <=32'h0021FFFA;
14'd11937:data <=32'h0022FFF5;14'd11938:data <=32'h0022FFEF;14'd11939:data <=32'h0020FFEA;
14'd11940:data <=32'h001CFFE5;14'd11941:data <=32'h0017FFE2;14'd11942:data <=32'h0012FFE1;
14'd11943:data <=32'h000DFFE2;14'd11944:data <=32'h000AFFE5;14'd11945:data <=32'h000AFFE8;
14'd11946:data <=32'h000BFFEA;14'd11947:data <=32'h000FFFEA;14'd11948:data <=32'h0012FFE7;
14'd11949:data <=32'h0014FFE2;14'd11950:data <=32'h0014FFDB;14'd11951:data <=32'h0011FFD3;
14'd11952:data <=32'h000BFFCD;14'd11953:data <=32'h0003FFC9;14'd11954:data <=32'hFFFBFFC7;
14'd11955:data <=32'hFFF3FFC7;14'd11956:data <=32'hFFECFFC9;14'd11957:data <=32'hFFE7FFCA;
14'd11958:data <=32'hFFE1FFCD;14'd11959:data <=32'hFFDBFFCF;14'd11960:data <=32'hFFD5FFD1;
14'd11961:data <=32'hFFCFFFD4;14'd11962:data <=32'hFFC9FFD9;14'd11963:data <=32'hFFC4FFDE;
14'd11964:data <=32'hFFBFFFE4;14'd11965:data <=32'hFFBBFFEA;14'd11966:data <=32'hFFB8FFEF;
14'd11967:data <=32'hFFB3FFF5;14'd11968:data <=32'hFFA5002E;14'd11969:data <=32'hFFAA003A;
14'd11970:data <=32'hFFB2003B;14'd11971:data <=32'hFFA30005;14'd11972:data <=32'hFF8B0002;
14'd11973:data <=32'hFF87001B;14'd11974:data <=32'hFF8A0034;14'd11975:data <=32'hFF95004E;
14'd11976:data <=32'hFFA60063;14'd11977:data <=32'hFFBB0073;14'd11978:data <=32'hFFD3007D;
14'd11979:data <=32'hFFED0080;14'd11980:data <=32'h0005007F;14'd11981:data <=32'h001D0079;
14'd11982:data <=32'h0032006D;14'd11983:data <=32'h0044005D;14'd11984:data <=32'h00510049;
14'd11985:data <=32'h00590033;14'd11986:data <=32'h0059001C;14'd11987:data <=32'h00540007;
14'd11988:data <=32'h0049FFF6;14'd11989:data <=32'h003AFFEB;14'd11990:data <=32'h002BFFE6;
14'd11991:data <=32'h001DFFE5;14'd11992:data <=32'h0012FFE9;14'd11993:data <=32'h000BFFEE;
14'd11994:data <=32'h0006FFF4;14'd11995:data <=32'h0004FFFA;14'd11996:data <=32'h0002FFFE;
14'd11997:data <=32'h00020003;14'd11998:data <=32'h00030007;14'd11999:data <=32'h0004000C;
14'd12000:data <=32'h00070010;14'd12001:data <=32'h000C0014;14'd12002:data <=32'h00120016;
14'd12003:data <=32'h00180016;14'd12004:data <=32'h001E0014;14'd12005:data <=32'h00240011;
14'd12006:data <=32'h0029000D;14'd12007:data <=32'h002C0008;14'd12008:data <=32'h00300003;
14'd12009:data <=32'h0033FFFD;14'd12010:data <=32'h0036FFF7;14'd12011:data <=32'h0038FFEE;
14'd12012:data <=32'h0039FFE5;14'd12013:data <=32'h0037FFDA;14'd12014:data <=32'h0032FFCF;
14'd12015:data <=32'h0029FFC4;14'd12016:data <=32'h001EFFBD;14'd12017:data <=32'h0010FFBA;
14'd12018:data <=32'h0003FFBB;14'd12019:data <=32'hFFF7FFC0;14'd12020:data <=32'hFFEFFFC8;
14'd12021:data <=32'hFFEBFFD0;14'd12022:data <=32'hFFE9FFD8;14'd12023:data <=32'hFFEBFFDE;
14'd12024:data <=32'hFFEDFFE1;14'd12025:data <=32'hFFF0FFE3;14'd12026:data <=32'hFFF3FFE2;
14'd12027:data <=32'hFFF5FFE0;14'd12028:data <=32'hFFF6FFDC;14'd12029:data <=32'hFFF6FFD6;
14'd12030:data <=32'hFFF3FFCF;14'd12031:data <=32'hFFECFFC7;14'd12032:data <=32'hFFC2FFD3;
14'd12033:data <=32'hFFB7FFD5;14'd12034:data <=32'hFFB6FFDC;14'd12035:data <=32'hFFD5FFD0;
14'd12036:data <=32'hFFB5FFC0;14'd12037:data <=32'hFFA4FFCD;14'd12038:data <=32'hFF98FFDF;
14'd12039:data <=32'hFF91FFF4;14'd12040:data <=32'hFF910009;14'd12041:data <=32'hFF96001D;
14'd12042:data <=32'hFF9E002F;14'd12043:data <=32'hFFA9003E;14'd12044:data <=32'hFFB6004A;
14'd12045:data <=32'hFFC50053;14'd12046:data <=32'hFFD5005A;14'd12047:data <=32'hFFE6005D;
14'd12048:data <=32'hFFF7005B;14'd12049:data <=32'h00070056;14'd12050:data <=32'h0014004D;
14'd12051:data <=32'h001E0042;14'd12052:data <=32'h00230037;14'd12053:data <=32'h0025002D;
14'd12054:data <=32'h00250024;14'd12055:data <=32'h0025001E;14'd12056:data <=32'h00240019;
14'd12057:data <=32'h00240014;14'd12058:data <=32'h0024000E;14'd12059:data <=32'h00230008;
14'd12060:data <=32'h00200001;14'd12061:data <=32'h001BFFFB;14'd12062:data <=32'h0014FFF7;
14'd12063:data <=32'h000BFFF6;14'd12064:data <=32'h0003FFF8;14'd12065:data <=32'hFFFCFFFD;
14'd12066:data <=32'hFFF70004;14'd12067:data <=32'hFFF5000D;14'd12068:data <=32'hFFF50016;
14'd12069:data <=32'hFFF9001F;14'd12070:data <=32'hFFFF0026;14'd12071:data <=32'h0007002C;
14'd12072:data <=32'h00110031;14'd12073:data <=32'h001E0033;14'd12074:data <=32'h002B0032;
14'd12075:data <=32'h003A002D;14'd12076:data <=32'h00470024;14'd12077:data <=32'h00520016;
14'd12078:data <=32'h00580005;14'd12079:data <=32'h0059FFF2;14'd12080:data <=32'h0055FFDF;
14'd12081:data <=32'h004BFFD0;14'd12082:data <=32'h003EFFC4;14'd12083:data <=32'h002FFFBE;
14'd12084:data <=32'h0021FFBC;14'd12085:data <=32'h0016FFBD;14'd12086:data <=32'h000CFFC1;
14'd12087:data <=32'h0006FFC6;14'd12088:data <=32'h0002FFCA;14'd12089:data <=32'hFFFFFFCE;
14'd12090:data <=32'hFFFDFFD1;14'd12091:data <=32'hFFFCFFD3;14'd12092:data <=32'hFFFCFFD4;
14'd12093:data <=32'hFFFEFFD3;14'd12094:data <=32'hFFFDFFD1;14'd12095:data <=32'hFFFDFFCC;
14'd12096:data <=32'h0011FFD8;14'd12097:data <=32'h000FFFC7;14'd12098:data <=32'h0004FFBF;
14'd12099:data <=32'hFFE4FFCF;14'd12100:data <=32'hFFCBFFBD;14'd12101:data <=32'hFFC0FFC7;
14'd12102:data <=32'hFFB8FFD3;14'd12103:data <=32'hFFB4FFE1;14'd12104:data <=32'hFFB4FFEF;
14'd12105:data <=32'hFFB8FFFB;14'd12106:data <=32'hFFBD0003;14'd12107:data <=32'hFFC30009;
14'd12108:data <=32'hFFC8000D;14'd12109:data <=32'hFFCC0010;14'd12110:data <=32'hFFCF0012;
14'd12111:data <=32'hFFD10015;14'd12112:data <=32'hFFD40018;14'd12113:data <=32'hFFD7001B;
14'd12114:data <=32'hFFD9001D;14'd12115:data <=32'hFFDB001F;14'd12116:data <=32'hFFDC0021;
14'd12117:data <=32'hFFDD0025;14'd12118:data <=32'hFFDF002A;14'd12119:data <=32'hFFE30030;
14'd12120:data <=32'hFFEA0037;14'd12121:data <=32'hFFF3003C;14'd12122:data <=32'h0000003D;
14'd12123:data <=32'h000C003A;14'd12124:data <=32'h00170033;14'd12125:data <=32'h001F0029;
14'd12126:data <=32'h0023001C;14'd12127:data <=32'h00220010;14'd12128:data <=32'h001D0006;
14'd12129:data <=32'h0016FFFF;14'd12130:data <=32'h000DFFFB;14'd12131:data <=32'h0004FFFB;
14'd12132:data <=32'hFFFCFFFD;14'd12133:data <=32'hFFF40001;14'd12134:data <=32'hFFEF0009;
14'd12135:data <=32'hFFEC0011;14'd12136:data <=32'hFFEB001B;14'd12137:data <=32'hFFED0026;
14'd12138:data <=32'hFFF30031;14'd12139:data <=32'hFFFD003A;14'd12140:data <=32'h000A0040;
14'd12141:data <=32'h00180041;14'd12142:data <=32'h0027003F;14'd12143:data <=32'h00350038;
14'd12144:data <=32'h003E002E;14'd12145:data <=32'h00450023;14'd12146:data <=32'h00490018;
14'd12147:data <=32'h004B000E;14'd12148:data <=32'h004B0005;14'd12149:data <=32'h004BFFFD;
14'd12150:data <=32'h004CFFF6;14'd12151:data <=32'h004DFFED;14'd12152:data <=32'h004DFFE3;
14'd12153:data <=32'h004BFFD8;14'd12154:data <=32'h0047FFCD;14'd12155:data <=32'h0041FFC1;
14'd12156:data <=32'h0038FFB8;14'd12157:data <=32'h002EFFB0;14'd12158:data <=32'h0023FFA9;
14'd12159:data <=32'h0017FFA4;14'd12160:data <=32'h0016FFFD;14'd12161:data <=32'h0024FFF1;
14'd12162:data <=32'h0029FFDA;14'd12163:data <=32'hFFFCFFA0;14'd12164:data <=32'hFFDAFF90;
14'd12165:data <=32'hFFC6FF9D;14'd12166:data <=32'hFFB7FFAF;14'd12167:data <=32'hFFAEFFC5;
14'd12168:data <=32'hFFACFFDA;14'd12169:data <=32'hFFB1FFEE;14'd12170:data <=32'hFFBBFFFC;
14'd12171:data <=32'hFFC60006;14'd12172:data <=32'hFFD1000A;14'd12173:data <=32'hFFDC000B;
14'd12174:data <=32'hFFE30009;14'd12175:data <=32'hFFE80005;14'd12176:data <=32'hFFEB0001;
14'd12177:data <=32'hFFEDFFFC;14'd12178:data <=32'hFFEBFFF8;14'd12179:data <=32'hFFE8FFF4;
14'd12180:data <=32'hFFE2FFF1;14'd12181:data <=32'hFFDAFFF2;14'd12182:data <=32'hFFD2FFF6;
14'd12183:data <=32'hFFCCFFFE;14'd12184:data <=32'hFFC80008;14'd12185:data <=32'hFFC90014;
14'd12186:data <=32'hFFCE0020;14'd12187:data <=32'hFFD60029;14'd12188:data <=32'hFFE1002E;
14'd12189:data <=32'hFFEC002F;14'd12190:data <=32'hFFF5002D;14'd12191:data <=32'hFFFC0029;
14'd12192:data <=32'h00010024;14'd12193:data <=32'h0004001E;14'd12194:data <=32'h00050019;
14'd12195:data <=32'h00050015;14'd12196:data <=32'h00040012;14'd12197:data <=32'h0003000F;
14'd12198:data <=32'h0000000D;14'd12199:data <=32'hFFFD000C;14'd12200:data <=32'hFFFA000B;
14'd12201:data <=32'hFFF6000D;14'd12202:data <=32'hFFF20010;14'd12203:data <=32'hFFF00015;
14'd12204:data <=32'hFFEF001A;14'd12205:data <=32'hFFF10020;14'd12206:data <=32'hFFF30025;
14'd12207:data <=32'hFFF60029;14'd12208:data <=32'hFFFA002D;14'd12209:data <=32'hFFFD0031;
14'd12210:data <=32'h00010036;14'd12211:data <=32'h0006003C;14'd12212:data <=32'h000D0042;
14'd12213:data <=32'h00180049;14'd12214:data <=32'h0027004D;14'd12215:data <=32'h0039004D;
14'd12216:data <=32'h004C0047;14'd12217:data <=32'h005F003D;14'd12218:data <=32'h006E002C;
14'd12219:data <=32'h007A0017;14'd12220:data <=32'h00810000;14'd12221:data <=32'h0081FFE7;
14'd12222:data <=32'h007DFFCF;14'd12223:data <=32'h0073FFB8;14'd12224:data <=32'h0025FFF2;
14'd12225:data <=32'h0031FFEC;14'd12226:data <=32'h0042FFE0;14'd12227:data <=32'h005EFFA9;
14'd12228:data <=32'h003AFF83;14'd12229:data <=32'h001EFF80;14'd12230:data <=32'h0003FF84;
14'd12231:data <=32'hFFEBFF8E;14'd12232:data <=32'hFFD9FF9D;14'd12233:data <=32'hFFCEFFAF;
14'd12234:data <=32'hFFC9FFC1;14'd12235:data <=32'hFFC9FFCF;14'd12236:data <=32'hFFCBFFDC;
14'd12237:data <=32'hFFCFFFE5;14'd12238:data <=32'hFFD3FFEC;14'd12239:data <=32'hFFD7FFF1;
14'd12240:data <=32'hFFDBFFF5;14'd12241:data <=32'hFFDFFFF7;14'd12242:data <=32'hFFE3FFF8;
14'd12243:data <=32'hFFE7FFF8;14'd12244:data <=32'hFFE8FFF6;14'd12245:data <=32'hFFE8FFF3;
14'd12246:data <=32'hFFE6FFF2;14'd12247:data <=32'hFFE3FFF3;14'd12248:data <=32'hFFDFFFF6;
14'd12249:data <=32'hFFDDFFFA;14'd12250:data <=32'hFFDDFFFE;14'd12251:data <=32'hFFDF0003;
14'd12252:data <=32'hFFE20005;14'd12253:data <=32'hFFE50006;14'd12254:data <=32'hFFE70005;
14'd12255:data <=32'hFFE70003;14'd12256:data <=32'hFFE50003;14'd12257:data <=32'hFFE20003;
14'd12258:data <=32'hFFDF0006;14'd12259:data <=32'hFFDE000B;14'd12260:data <=32'hFFDE0010;
14'd12261:data <=32'hFFE00015;14'd12262:data <=32'hFFE4001A;14'd12263:data <=32'hFFE9001C;
14'd12264:data <=32'hFFED001D;14'd12265:data <=32'hFFF1001D;14'd12266:data <=32'hFFF5001C;
14'd12267:data <=32'hFFF7001A;14'd12268:data <=32'hFFF90018;14'd12269:data <=32'hFFFA0015;
14'd12270:data <=32'hFFF90012;14'd12271:data <=32'hFFF7000F;14'd12272:data <=32'hFFF3000D;
14'd12273:data <=32'hFFED000D;14'd12274:data <=32'hFFE50011;14'd12275:data <=32'hFFDD0019;
14'd12276:data <=32'hFFD80024;14'd12277:data <=32'hFFD70034;14'd12278:data <=32'hFFDC0045;
14'd12279:data <=32'hFFE80055;14'd12280:data <=32'hFFF90062;14'd12281:data <=32'h000F006A;
14'd12282:data <=32'h0026006C;14'd12283:data <=32'h003D0067;14'd12284:data <=32'h0053005C;
14'd12285:data <=32'h0066004D;14'd12286:data <=32'h0074003A;14'd12287:data <=32'h007F0024;
14'd12288:data <=32'h00540024;14'd12289:data <=32'h00660019;14'd12290:data <=32'h00730011;
14'd12291:data <=32'h007A0013;14'd12292:data <=32'h006BFFE6;14'd12293:data <=32'h0062FFD6;
14'd12294:data <=32'h0055FFCA;14'd12295:data <=32'h0048FFC1;14'd12296:data <=32'h003BFFBD;
14'd12297:data <=32'h0031FFBB;14'd12298:data <=32'h0028FFBA;14'd12299:data <=32'h0021FFB8;
14'd12300:data <=32'h001AFFB6;14'd12301:data <=32'h0011FFB4;14'd12302:data <=32'h0007FFB2;
14'd12303:data <=32'hFFFBFFB2;14'd12304:data <=32'hFFF0FFB4;14'd12305:data <=32'hFFE5FFBB;
14'd12306:data <=32'hFFDCFFC2;14'd12307:data <=32'hFFD6FFCC;14'd12308:data <=32'hFFD1FFD6;
14'd12309:data <=32'hFFCFFFDF;14'd12310:data <=32'hFFCEFFE9;14'd12311:data <=32'hFFCFFFF2;
14'd12312:data <=32'hFFD2FFFB;14'd12313:data <=32'hFFD70004;14'd12314:data <=32'hFFDE000A;
14'd12315:data <=32'hFFE8000E;14'd12316:data <=32'hFFF3000E;14'd12317:data <=32'hFFFC000A;
14'd12318:data <=32'h00030002;14'd12319:data <=32'h0006FFF9;14'd12320:data <=32'h0004FFEE;
14'd12321:data <=32'hFFFEFFE6;14'd12322:data <=32'hFFF5FFE1;14'd12323:data <=32'hFFECFFDF;
14'd12324:data <=32'hFFE2FFE2;14'd12325:data <=32'hFFDAFFE7;14'd12326:data <=32'hFFD5FFED;
14'd12327:data <=32'hFFD1FFF5;14'd12328:data <=32'hFFD0FFFC;14'd12329:data <=32'hFFD00003;
14'd12330:data <=32'hFFD20009;14'd12331:data <=32'hFFD5000F;14'd12332:data <=32'hFFD80013;
14'd12333:data <=32'hFFDC0017;14'd12334:data <=32'hFFE10018;14'd12335:data <=32'hFFE50018;
14'd12336:data <=32'hFFE70016;14'd12337:data <=32'hFFE60014;14'd12338:data <=32'hFFE40013;
14'd12339:data <=32'hFFDF0013;14'd12340:data <=32'hFFDA0017;14'd12341:data <=32'hFFD6001F;
14'd12342:data <=32'hFFD4002A;14'd12343:data <=32'hFFD60037;14'd12344:data <=32'hFFDD0042;
14'd12345:data <=32'hFFE8004C;14'd12346:data <=32'hFFF50053;14'd12347:data <=32'h00030056;
14'd12348:data <=32'h00110056;14'd12349:data <=32'h001D0053;14'd12350:data <=32'h002A004D;
14'd12351:data <=32'h00340047;14'd12352:data <=32'h00200074;14'd12353:data <=32'h00400077;
14'd12354:data <=32'h0055006C;14'd12355:data <=32'h00360042;14'd12356:data <=32'h00300024;
14'd12357:data <=32'h00310021;14'd12358:data <=32'h0033001E;14'd12359:data <=32'h0035001C;
14'd12360:data <=32'h003A001B;14'd12361:data <=32'h0040001A;14'd12362:data <=32'h00490015;
14'd12363:data <=32'h0052000D;14'd12364:data <=32'h005AFFFF;14'd12365:data <=32'h005FFFEE;
14'd12366:data <=32'h005EFFDB;14'd12367:data <=32'h0056FFC8;14'd12368:data <=32'h004AFFB8;
14'd12369:data <=32'h003AFFAC;14'd12370:data <=32'h0028FFA4;14'd12371:data <=32'h0015FFA1;
14'd12372:data <=32'h0003FFA3;14'd12373:data <=32'hFFF2FFA8;14'd12374:data <=32'hFFE3FFB1;
14'd12375:data <=32'hFFD6FFBD;14'd12376:data <=32'hFFCCFFCB;14'd12377:data <=32'hFFC7FFDC;
14'd12378:data <=32'hFFC8FFED;14'd12379:data <=32'hFFCDFFFD;14'd12380:data <=32'hFFD70009;
14'd12381:data <=32'hFFE50011;14'd12382:data <=32'hFFF20013;14'd12383:data <=32'hFFFF0010;
14'd12384:data <=32'h00090009;14'd12385:data <=32'h000FFFFF;14'd12386:data <=32'h0011FFF6;
14'd12387:data <=32'h0010FFED;14'd12388:data <=32'h000CFFE6;14'd12389:data <=32'h0008FFE0;
14'd12390:data <=32'h0003FFDC;14'd12391:data <=32'hFFFDFFD8;14'd12392:data <=32'hFFF7FFD5;
14'd12393:data <=32'hFFF0FFD3;14'd12394:data <=32'hFFE8FFD2;14'd12395:data <=32'hFFE0FFD3;
14'd12396:data <=32'hFFD7FFD6;14'd12397:data <=32'hFFCFFFDA;14'd12398:data <=32'hFFC8FFE0;
14'd12399:data <=32'hFFC3FFE7;14'd12400:data <=32'hFFBEFFEF;14'd12401:data <=32'hFFBAFFF7;
14'd12402:data <=32'hFFB70000;14'd12403:data <=32'hFFB40009;14'd12404:data <=32'hFFB20015;
14'd12405:data <=32'hFFB20022;14'd12406:data <=32'hFFB60030;14'd12407:data <=32'hFFBD003E;
14'd12408:data <=32'hFFC9004A;14'd12409:data <=32'hFFD80053;14'd12410:data <=32'hFFE90057;
14'd12411:data <=32'hFFF90055;14'd12412:data <=32'h00080050;14'd12413:data <=32'h00120048;
14'd12414:data <=32'h0019003E;14'd12415:data <=32'h001D0036;14'd12416:data <=32'hFFCC005B;
14'd12417:data <=32'hFFDE0071;14'd12418:data <=32'hFFFA0077;14'd12419:data <=32'h001D0038;
14'd12420:data <=32'h0011001B;14'd12421:data <=32'h000C001A;14'd12422:data <=32'h0008001D;
14'd12423:data <=32'h00050023;14'd12424:data <=32'h0006002B;14'd12425:data <=32'h000B0034;
14'd12426:data <=32'h0015003C;14'd12427:data <=32'h00230040;14'd12428:data <=32'h0034003F;
14'd12429:data <=32'h00440037;14'd12430:data <=32'h0052002A;14'd12431:data <=32'h005B001A;
14'd12432:data <=32'h005F0007;14'd12433:data <=32'h005EFFF5;14'd12434:data <=32'h0058FFE4;
14'd12435:data <=32'h0050FFD6;14'd12436:data <=32'h0045FFCA;14'd12437:data <=32'h0038FFC2;
14'd12438:data <=32'h002BFFBB;14'd12439:data <=32'h001CFFB8;14'd12440:data <=32'h000DFFB9;
14'd12441:data <=32'hFFFEFFBE;14'd12442:data <=32'hFFF3FFC6;14'd12443:data <=32'hFFEBFFD0;
14'd12444:data <=32'hFFE6FFDC;14'd12445:data <=32'hFFE6FFE7;14'd12446:data <=32'hFFE8FFF0;
14'd12447:data <=32'hFFEDFFF7;14'd12448:data <=32'hFFF2FFFB;14'd12449:data <=32'hFFF7FFFD;
14'd12450:data <=32'hFFFBFFFE;14'd12451:data <=32'hFFFF0000;14'd12452:data <=32'h00030000;
14'd12453:data <=32'h00080000;14'd12454:data <=32'h000EFFFF;14'd12455:data <=32'h0015FFFC;
14'd12456:data <=32'h001CFFF5;14'd12457:data <=32'h0021FFEC;14'd12458:data <=32'h0022FFE0;
14'd12459:data <=32'h0021FFD3;14'd12460:data <=32'h001AFFC7;14'd12461:data <=32'h0011FFBC;
14'd12462:data <=32'h0004FFB3;14'd12463:data <=32'hFFF5FFAD;14'd12464:data <=32'hFFE4FFAA;
14'd12465:data <=32'hFFD3FFAB;14'd12466:data <=32'hFFC0FFB0;14'd12467:data <=32'hFFAEFFB9;
14'd12468:data <=32'hFF9EFFC7;14'd12469:data <=32'hFF90FFDA;14'd12470:data <=32'hFF88FFF1;
14'd12471:data <=32'hFF85000A;14'd12472:data <=32'hFF8A0023;14'd12473:data <=32'hFF96003A;
14'd12474:data <=32'hFFA7004C;14'd12475:data <=32'hFFBC0057;14'd12476:data <=32'hFFD1005C;
14'd12477:data <=32'hFFE4005B;14'd12478:data <=32'hFFF50055;14'd12479:data <=32'h0001004D;
14'd12480:data <=32'hFFCD0029;14'd12481:data <=32'hFFCD0038;14'd12482:data <=32'hFFD7004B;
14'd12483:data <=32'h00010058;14'd12484:data <=32'hFFFF0039;14'd12485:data <=32'h00010035;
14'd12486:data <=32'h00020032;14'd12487:data <=32'h00030031;14'd12488:data <=32'h00030032;
14'd12489:data <=32'h00050035;14'd12490:data <=32'h000A0039;14'd12491:data <=32'h0011003C;
14'd12492:data <=32'h001C003D;14'd12493:data <=32'h00270039;14'd12494:data <=32'h00300033;
14'd12495:data <=32'h00370029;14'd12496:data <=32'h003B001E;14'd12497:data <=32'h003B0014;
14'd12498:data <=32'h0039000B;14'd12499:data <=32'h00360004;14'd12500:data <=32'h00330000;
14'd12501:data <=32'h0030FFFB;14'd12502:data <=32'h002EFFF8;14'd12503:data <=32'h002CFFF4;
14'd12504:data <=32'h0028FFF0;14'd12505:data <=32'h0025FFED;14'd12506:data <=32'h0020FFEB;
14'd12507:data <=32'h001DFFEA;14'd12508:data <=32'h001AFFE9;14'd12509:data <=32'h0017FFE9;
14'd12510:data <=32'h0016FFE8;14'd12511:data <=32'h0014FFE7;14'd12512:data <=32'h0011FFE5;
14'd12513:data <=32'h000CFFE3;14'd12514:data <=32'h0006FFE3;14'd12515:data <=32'h0001FFE6;
14'd12516:data <=32'hFFFCFFEB;14'd12517:data <=32'hFFF9FFF2;14'd12518:data <=32'hFFFAFFFB;
14'd12519:data <=32'hFFFF0003;14'd12520:data <=32'h00070009;14'd12521:data <=32'h0012000A;
14'd12522:data <=32'h001E0007;14'd12523:data <=32'h00280001;14'd12524:data <=32'h0030FFF6;
14'd12525:data <=32'h0034FFE9;14'd12526:data <=32'h0035FFDA;14'd12527:data <=32'h0032FFCB;
14'd12528:data <=32'h002BFFBD;14'd12529:data <=32'h0021FFAF;14'd12530:data <=32'h0013FFA4;
14'd12531:data <=32'h0001FF9C;14'd12532:data <=32'hFFECFF97;14'd12533:data <=32'hFFD7FF99;
14'd12534:data <=32'hFFC1FFA1;14'd12535:data <=32'hFFAEFFAE;14'd12536:data <=32'hFFA0FFC0;
14'd12537:data <=32'hFF97FFD4;14'd12538:data <=32'hFF95FFE9;14'd12539:data <=32'hFF97FFFC;
14'd12540:data <=32'hFF9D000B;14'd12541:data <=32'hFFA40017;14'd12542:data <=32'hFFAC0021;
14'd12543:data <=32'hFFB30028;14'd12544:data <=32'hFFC5002C;14'd12545:data <=32'hFFC80032;
14'd12546:data <=32'hFFC6003A;14'd12547:data <=32'hFFA8003C;14'd12548:data <=32'hFFA90030;
14'd12549:data <=32'hFFB0003C;14'd12550:data <=32'hFFB90047;14'd12551:data <=32'hFFC50051;
14'd12552:data <=32'hFFD20059;14'd12553:data <=32'hFFDF0060;14'd12554:data <=32'hFFF00064;
14'd12555:data <=32'h00010064;14'd12556:data <=32'h00140061;14'd12557:data <=32'h00260058;
14'd12558:data <=32'h0034004B;14'd12559:data <=32'h003E003A;14'd12560:data <=32'h00410028;
14'd12561:data <=32'h003F0017;14'd12562:data <=32'h00380009;14'd12563:data <=32'h002FFFFF;
14'd12564:data <=32'h0024FFFA;14'd12565:data <=32'h001BFFFA;14'd12566:data <=32'h0013FFFC;
14'd12567:data <=32'h000EFFFE;14'd12568:data <=32'h000B0003;14'd12569:data <=32'h00090007;
14'd12570:data <=32'h000A000C;14'd12571:data <=32'h000C0010;14'd12572:data <=32'h000F0014;
14'd12573:data <=32'h00150015;14'd12574:data <=32'h001C0015;14'd12575:data <=32'h00220011;
14'd12576:data <=32'h0027000C;14'd12577:data <=32'h002A0003;14'd12578:data <=32'h0029FFFB;
14'd12579:data <=32'h0025FFF4;14'd12580:data <=32'h001FFFF0;14'd12581:data <=32'h0018FFEF;
14'd12582:data <=32'h0013FFF1;14'd12583:data <=32'h000FFFF5;14'd12584:data <=32'h0010FFFA;
14'd12585:data <=32'h0012FFFE;14'd12586:data <=32'h00160000;14'd12587:data <=32'h001CFFFF;
14'd12588:data <=32'h0021FFFD;14'd12589:data <=32'h0025FFF9;14'd12590:data <=32'h0028FFF3;
14'd12591:data <=32'h002AFFED;14'd12592:data <=32'h002BFFE6;14'd12593:data <=32'h002BFFDF;
14'd12594:data <=32'h002AFFD6;14'd12595:data <=32'h0027FFCE;14'd12596:data <=32'h0021FFC6;
14'd12597:data <=32'h0019FFBE;14'd12598:data <=32'h000FFFB9;14'd12599:data <=32'h0005FFB6;
14'd12600:data <=32'hFFFBFFB7;14'd12601:data <=32'hFFF2FFB8;14'd12602:data <=32'hFFEBFFBA;
14'd12603:data <=32'hFFE5FFBC;14'd12604:data <=32'hFFDEFFBC;14'd12605:data <=32'hFFD7FFBC;
14'd12606:data <=32'hFFCEFFBC;14'd12607:data <=32'hFFC1FFBD;14'd12608:data <=32'hFFA5FFF6;
14'd12609:data <=32'hFFA30001;14'd12610:data <=32'hFFA60004;14'd12611:data <=32'hFFA5FFCE;
14'd12612:data <=32'hFF91FFC4;14'd12613:data <=32'hFF85FFD9;14'd12614:data <=32'hFF7DFFF0;
14'd12615:data <=32'hFF7B0009;14'd12616:data <=32'hFF7E0022;14'd12617:data <=32'hFF87003A;
14'd12618:data <=32'hFF950051;14'd12619:data <=32'hFFA90064;14'd12620:data <=32'hFFC10071;
14'd12621:data <=32'hFFDC0077;14'd12622:data <=32'hFFF70075;14'd12623:data <=32'h0010006C;
14'd12624:data <=32'h0023005D;14'd12625:data <=32'h0030004A;14'd12626:data <=32'h00350037;
14'd12627:data <=32'h00360025;14'd12628:data <=32'h00310017;14'd12629:data <=32'h002B000C;
14'd12630:data <=32'h00230004;14'd12631:data <=32'h001BFFFF;14'd12632:data <=32'h0014FFFD;
14'd12633:data <=32'h000CFFFC;14'd12634:data <=32'h0005FFFE;14'd12635:data <=32'hFFFF0001;
14'd12636:data <=32'hFFFB0007;14'd12637:data <=32'hFFF9000E;14'd12638:data <=32'hFFFA0014;
14'd12639:data <=32'hFFFE001A;14'd12640:data <=32'h0003001E;14'd12641:data <=32'h0009001F;
14'd12642:data <=32'h000E001F;14'd12643:data <=32'h0011001D;14'd12644:data <=32'h0014001C;
14'd12645:data <=32'h0016001C;14'd12646:data <=32'h0019001B;14'd12647:data <=32'h001D001C;
14'd12648:data <=32'h0023001C;14'd12649:data <=32'h0029001A;14'd12650:data <=32'h00310016;
14'd12651:data <=32'h0036000E;14'd12652:data <=32'h003A0006;14'd12653:data <=32'h003CFFFC;
14'd12654:data <=32'h0039FFF2;14'd12655:data <=32'h0035FFE9;14'd12656:data <=32'h0030FFE3;
14'd12657:data <=32'h0029FFDF;14'd12658:data <=32'h0023FFDD;14'd12659:data <=32'h001EFFDC;
14'd12660:data <=32'h0019FFDC;14'd12661:data <=32'h0016FFDD;14'd12662:data <=32'h0012FFDE;
14'd12663:data <=32'h0011FFE1;14'd12664:data <=32'h0011FFE3;14'd12665:data <=32'h0014FFE5;
14'd12666:data <=32'h0018FFE4;14'd12667:data <=32'h001EFFE1;14'd12668:data <=32'h0023FFD8;
14'd12669:data <=32'h0026FFCC;14'd12670:data <=32'h0024FFBD;14'd12671:data <=32'h001CFFAD;
14'd12672:data <=32'hFFE6FFB3;14'd12673:data <=32'hFFDAFFAF;14'd12674:data <=32'hFFD6FFB4;
14'd12675:data <=32'hFFF9FFAE;14'd12676:data <=32'hFFE1FF93;14'd12677:data <=32'hFFCBFF98;
14'd12678:data <=32'hFFB8FFA2;14'd12679:data <=32'hFFA7FFAF;14'd12680:data <=32'hFF9AFFC0;
14'd12681:data <=32'hFF8FFFD4;14'd12682:data <=32'hFF89FFEA;14'd12683:data <=32'hFF890002;
14'd12684:data <=32'hFF8F0019;14'd12685:data <=32'hFF9A002C;14'd12686:data <=32'hFFAA003C;
14'd12687:data <=32'hFFBC0045;14'd12688:data <=32'hFFCE0049;14'd12689:data <=32'hFFDD0048;
14'd12690:data <=32'hFFEA0045;14'd12691:data <=32'hFFF40040;14'd12692:data <=32'hFFFB003B;
14'd12693:data <=32'h00010037;14'd12694:data <=32'h00070033;14'd12695:data <=32'h000C002D;
14'd12696:data <=32'h00110027;14'd12697:data <=32'h00150020;14'd12698:data <=32'h00160018;
14'd12699:data <=32'h00150011;14'd12700:data <=32'h0012000A;14'd12701:data <=32'h000D0006;
14'd12702:data <=32'h00080003;14'd12703:data <=32'h00030002;14'd12704:data <=32'hFFFE0002;
14'd12705:data <=32'hFFF90003;14'd12706:data <=32'hFFF40006;14'd12707:data <=32'hFFEF000A;
14'd12708:data <=32'hFFEB0010;14'd12709:data <=32'hFFE80019;14'd12710:data <=32'hFFE80023;
14'd12711:data <=32'hFFEC002E;14'd12712:data <=32'hFFF40039;14'd12713:data <=32'h00000042;
14'd12714:data <=32'h000F0046;14'd12715:data <=32'h00200045;14'd12716:data <=32'h002F003F;
14'd12717:data <=32'h003C0035;14'd12718:data <=32'h00460028;14'd12719:data <=32'h004B001A;
14'd12720:data <=32'h004C000C;14'd12721:data <=32'h0049FFFF;14'd12722:data <=32'h0044FFF4;
14'd12723:data <=32'h003EFFEC;14'd12724:data <=32'h0037FFE6;14'd12725:data <=32'h0030FFE1;
14'd12726:data <=32'h0028FFE0;14'd12727:data <=32'h0021FFE0;14'd12728:data <=32'h001CFFE3;
14'd12729:data <=32'h0019FFE7;14'd12730:data <=32'h001AFFEC;14'd12731:data <=32'h001FFFEF;
14'd12732:data <=32'h0026FFEE;14'd12733:data <=32'h002DFFE9;14'd12734:data <=32'h0033FFDF;
14'd12735:data <=32'h0035FFD2;14'd12736:data <=32'h0036FFE0;14'd12737:data <=32'h003AFFCD;
14'd12738:data <=32'h0033FFC1;14'd12739:data <=32'h0014FFC8;14'd12740:data <=32'h0006FFAC;
14'd12741:data <=32'hFFF9FFAD;14'd12742:data <=32'hFFEEFFB0;14'd12743:data <=32'hFFE4FFB6;
14'd12744:data <=32'hFFDCFFBC;14'd12745:data <=32'hFFD4FFC2;14'd12746:data <=32'hFFCDFFCA;
14'd12747:data <=32'hFFC8FFD3;14'd12748:data <=32'hFFC5FFDC;14'd12749:data <=32'hFFC5FFE5;
14'd12750:data <=32'hFFC6FFED;14'd12751:data <=32'hFFC8FFF2;14'd12752:data <=32'hFFCBFFF6;
14'd12753:data <=32'hFFCBFFF8;14'd12754:data <=32'hFFCAFFFA;14'd12755:data <=32'hFFC7FFFE;
14'd12756:data <=32'hFFC40005;14'd12757:data <=32'hFFC2000E;14'd12758:data <=32'hFFC40018;
14'd12759:data <=32'hFFC80023;14'd12760:data <=32'hFFD1002C;14'd12761:data <=32'hFFDC0033;
14'd12762:data <=32'hFFE80035;14'd12763:data <=32'hFFF40034;14'd12764:data <=32'hFFFE0030;
14'd12765:data <=32'h0006002A;14'd12766:data <=32'h000C0023;14'd12767:data <=32'h0010001A;
14'd12768:data <=32'h00110011;14'd12769:data <=32'h000F0008;14'd12770:data <=32'h000BFFFF;
14'd12771:data <=32'h0003FFF8;14'd12772:data <=32'hFFF9FFF4;14'd12773:data <=32'hFFEEFFF5;
14'd12774:data <=32'hFFE2FFFA;14'd12775:data <=32'hFFD80003;14'd12776:data <=32'hFFD30010;
14'd12777:data <=32'hFFD2001F;14'd12778:data <=32'hFFD6002D;14'd12779:data <=32'hFFDE0039;
14'd12780:data <=32'hFFEA0042;14'd12781:data <=32'hFFF70047;14'd12782:data <=32'h00030048;
14'd12783:data <=32'h000F0047;14'd12784:data <=32'h00190044;14'd12785:data <=32'h00220040;
14'd12786:data <=32'h002B003C;14'd12787:data <=32'h00320036;14'd12788:data <=32'h00390030;
14'd12789:data <=32'h003F0029;14'd12790:data <=32'h00440021;14'd12791:data <=32'h00470018;
14'd12792:data <=32'h00490010;14'd12793:data <=32'h004A0008;14'd12794:data <=32'h004B0001;
14'd12795:data <=32'h004DFFFA;14'd12796:data <=32'h004FFFF1;14'd12797:data <=32'h0050FFE7;
14'd12798:data <=32'h004FFFDB;14'd12799:data <=32'h004CFFCD;14'd12800:data <=32'h00270019;
14'd12801:data <=32'h003C0011;14'd12802:data <=32'h0048FFFC;14'd12803:data <=32'h002EFFBA;
14'd12804:data <=32'h0019FF9D;14'd12805:data <=32'h0006FFA2;14'd12806:data <=32'hFFF7FFAB;
14'd12807:data <=32'hFFEBFFB6;14'd12808:data <=32'hFFE4FFC2;14'd12809:data <=32'hFFE1FFCD;
14'd12810:data <=32'hFFE0FFD7;14'd12811:data <=32'hFFE1FFE0;14'd12812:data <=32'hFFE4FFE7;
14'd12813:data <=32'hFFEAFFEC;14'd12814:data <=32'hFFF0FFEE;14'd12815:data <=32'hFFF6FFED;
14'd12816:data <=32'hFFFBFFE8;14'd12817:data <=32'hFFFCFFE1;14'd12818:data <=32'hFFF8FFD9;
14'd12819:data <=32'hFFF0FFD2;14'd12820:data <=32'hFFE6FFCF;14'd12821:data <=32'hFFD9FFD1;
14'd12822:data <=32'hFFCEFFD7;14'd12823:data <=32'hFFC5FFE2;14'd12824:data <=32'hFFC0FFEE;
14'd12825:data <=32'hFFBFFFFB;14'd12826:data <=32'hFFC20007;14'd12827:data <=32'hFFC80011;
14'd12828:data <=32'hFFCF0019;14'd12829:data <=32'hFFD7001E;14'd12830:data <=32'hFFDF0021;
14'd12831:data <=32'hFFE70022;14'd12832:data <=32'hFFF00022;14'd12833:data <=32'hFFF8001E;
14'd12834:data <=32'hFFFE0019;14'd12835:data <=32'h00020012;14'd12836:data <=32'h0003000A;
14'd12837:data <=32'h00000002;14'd12838:data <=32'hFFFBFFFC;14'd12839:data <=32'hFFF4FFF9;
14'd12840:data <=32'hFFECFFFA;14'd12841:data <=32'hFFE6FFFD;14'd12842:data <=32'hFFE10002;
14'd12843:data <=32'hFFDE0007;14'd12844:data <=32'hFFDD000C;14'd12845:data <=32'hFFDB0011;
14'd12846:data <=32'hFFDA0015;14'd12847:data <=32'hFFD8001A;14'd12848:data <=32'hFFD60021;
14'd12849:data <=32'hFFD5002A;14'd12850:data <=32'hFFD60034;14'd12851:data <=32'hFFDA0041;
14'd12852:data <=32'hFFE2004D;14'd12853:data <=32'hFFED0058;14'd12854:data <=32'hFFFC0060;
14'd12855:data <=32'h000D0065;14'd12856:data <=32'h001F0066;14'd12857:data <=32'h00320064;
14'd12858:data <=32'h0045005E;14'd12859:data <=32'h00570054;14'd12860:data <=32'h00690046;
14'd12861:data <=32'h00780034;14'd12862:data <=32'h0083001D;14'd12863:data <=32'h00880002;
14'd12864:data <=32'h00230018;14'd12865:data <=32'h00320019;14'd12866:data <=32'h00480015;
14'd12867:data <=32'h0077FFE5;14'd12868:data <=32'h0065FFB7;14'd12869:data <=32'h004FFFAC;
14'd12870:data <=32'h003AFFA7;14'd12871:data <=32'h0026FFA7;14'd12872:data <=32'h0015FFAC;
14'd12873:data <=32'h0007FFB2;14'd12874:data <=32'hFFFDFFBB;14'd12875:data <=32'hFFF5FFC4;
14'd12876:data <=32'hFFF0FFCE;14'd12877:data <=32'hFFEFFFD8;14'd12878:data <=32'hFFF0FFE0;
14'd12879:data <=32'hFFF4FFE6;14'd12880:data <=32'hFFFAFFE9;14'd12881:data <=32'hFFFFFFE8;
14'd12882:data <=32'h0002FFE4;14'd12883:data <=32'h0002FFDF;14'd12884:data <=32'hFFFFFFDA;
14'd12885:data <=32'hFFF8FFD6;14'd12886:data <=32'hFFF1FFD7;14'd12887:data <=32'hFFEAFFD9;
14'd12888:data <=32'hFFE6FFDE;14'd12889:data <=32'hFFE3FFE3;14'd12890:data <=32'hFFE2FFE7;
14'd12891:data <=32'hFFE2FFEB;14'd12892:data <=32'hFFE2FFEE;14'd12893:data <=32'hFFE1FFEF;
14'd12894:data <=32'hFFE0FFF1;14'd12895:data <=32'hFFE0FFF4;14'd12896:data <=32'hFFDFFFF7;
14'd12897:data <=32'hFFDFFFFB;14'd12898:data <=32'hFFE0FFFE;14'd12899:data <=32'hFFE20001;
14'd12900:data <=32'hFFE40002;14'd12901:data <=32'hFFE50003;14'd12902:data <=32'hFFE60004;
14'd12903:data <=32'hFFE70005;14'd12904:data <=32'hFFE80007;14'd12905:data <=32'hFFE90009;
14'd12906:data <=32'hFFEC000A;14'd12907:data <=32'hFFEF0009;14'd12908:data <=32'hFFF20006;
14'd12909:data <=32'hFFF30001;14'd12910:data <=32'hFFF2FFFB;14'd12911:data <=32'hFFECFFF5;
14'd12912:data <=32'hFFE3FFF1;14'd12913:data <=32'hFFD8FFF0;14'd12914:data <=32'hFFCAFFF5;
14'd12915:data <=32'hFFBFFFFF;14'd12916:data <=32'hFFB5000E;14'd12917:data <=32'hFFB1001F;
14'd12918:data <=32'hFFB10033;14'd12919:data <=32'hFFB70046;14'd12920:data <=32'hFFC10059;
14'd12921:data <=32'hFFCF0069;14'd12922:data <=32'hFFE20076;14'd12923:data <=32'hFFF80080;
14'd12924:data <=32'h00120084;14'd12925:data <=32'h002D0083;14'd12926:data <=32'h00480079;
14'd12927:data <=32'h00600069;14'd12928:data <=32'h0031004A;14'd12929:data <=32'h00450049;
14'd12930:data <=32'h00540049;14'd12931:data <=32'h00620050;14'd12932:data <=32'h00660023;
14'd12933:data <=32'h00640013;14'd12934:data <=32'h00600005;14'd12935:data <=32'h005BFFFB;
14'd12936:data <=32'h0056FFF0;14'd12937:data <=32'h0051FFE7;14'd12938:data <=32'h004CFFDE;
14'd12939:data <=32'h0045FFD6;14'd12940:data <=32'h003DFFCF;14'd12941:data <=32'h0033FFCA;
14'd12942:data <=32'h002BFFC7;14'd12943:data <=32'h0022FFC6;14'd12944:data <=32'h001BFFC5;
14'd12945:data <=32'h0014FFC4;14'd12946:data <=32'h000CFFC4;14'd12947:data <=32'h0004FFC3;
14'd12948:data <=32'hFFFBFFC5;14'd12949:data <=32'hFFF1FFCA;14'd12950:data <=32'hFFE9FFD1;
14'd12951:data <=32'hFFE3FFDB;14'd12952:data <=32'hFFE2FFE6;14'd12953:data <=32'hFFE4FFF0;
14'd12954:data <=32'hFFEAFFF8;14'd12955:data <=32'hFFF2FFFC;14'd12956:data <=32'hFFFAFFFD;
14'd12957:data <=32'h0001FFFA;14'd12958:data <=32'h0006FFF5;14'd12959:data <=32'h0007FFEF;
14'd12960:data <=32'h0007FFE9;14'd12961:data <=32'h0004FFE4;14'd12962:data <=32'h0000FFE0;
14'd12963:data <=32'hFFFBFFDD;14'd12964:data <=32'hFFF4FFDB;14'd12965:data <=32'hFFEEFFDB;
14'd12966:data <=32'hFFE7FFDC;14'd12967:data <=32'hFFE1FFE0;14'd12968:data <=32'hFFDBFFE5;
14'd12969:data <=32'hFFD8FFEC;14'd12970:data <=32'hFFD8FFF4;14'd12971:data <=32'hFFDAFFFB;
14'd12972:data <=32'hFFDFFFFF;14'd12973:data <=32'hFFE50000;14'd12974:data <=32'hFFE9FFFE;
14'd12975:data <=32'hFFECFFF9;14'd12976:data <=32'hFFEBFFF3;14'd12977:data <=32'hFFE5FFEE;
14'd12978:data <=32'hFFDDFFEB;14'd12979:data <=32'hFFD3FFEC;14'd12980:data <=32'hFFC9FFF0;
14'd12981:data <=32'hFFC0FFF9;14'd12982:data <=32'hFFBA0004;14'd12983:data <=32'hFFB60010;
14'd12984:data <=32'hFFB5001D;14'd12985:data <=32'hFFB6002B;14'd12986:data <=32'hFFBA0038;
14'd12987:data <=32'hFFC10046;14'd12988:data <=32'hFFCC0052;14'd12989:data <=32'hFFDA005D;
14'd12990:data <=32'hFFEA0064;14'd12991:data <=32'hFFFC0067;14'd12992:data <=32'hFFE5007B;
14'd12993:data <=32'hFFFE0088;14'd12994:data <=32'h00130088;14'd12995:data <=32'h0003005D;
14'd12996:data <=32'h00090041;14'd12997:data <=32'h000D0042;14'd12998:data <=32'h00110045;
14'd12999:data <=32'h00180049;14'd13000:data <=32'h0024004B;14'd13001:data <=32'h0031004A;
14'd13002:data <=32'h003F0045;14'd13003:data <=32'h004D003C;14'd13004:data <=32'h0059002E;
14'd13005:data <=32'h0060001F;14'd13006:data <=32'h0065000E;14'd13007:data <=32'h0066FFFD;
14'd13008:data <=32'h0064FFEB;14'd13009:data <=32'h005EFFDA;14'd13010:data <=32'h0054FFCA;
14'd13011:data <=32'h0046FFBC;14'd13012:data <=32'h0035FFB2;14'd13013:data <=32'h0021FFAC;
14'd13014:data <=32'h000CFFAD;14'd13015:data <=32'hFFF9FFB4;14'd13016:data <=32'hFFEAFFC1;
14'd13017:data <=32'hFFE1FFD0;14'd13018:data <=32'hFFDDFFE1;14'd13019:data <=32'hFFDFFFEF;
14'd13020:data <=32'hFFE6FFFC;14'd13021:data <=32'hFFEF0004;14'd13022:data <=32'hFFF80007;
14'd13023:data <=32'h00010008;14'd13024:data <=32'h000A0006;14'd13025:data <=32'h00110002;
14'd13026:data <=32'h0016FFFD;14'd13027:data <=32'h001AFFF6;14'd13028:data <=32'h001CFFEF;
14'd13029:data <=32'h001CFFE7;14'd13030:data <=32'h001AFFDE;14'd13031:data <=32'h0015FFD7;
14'd13032:data <=32'h000EFFD1;14'd13033:data <=32'h0006FFCD;14'd13034:data <=32'hFFFEFFCC;
14'd13035:data <=32'hFFF7FFCD;14'd13036:data <=32'hFFF1FFCE;14'd13037:data <=32'hFFEDFFCF;
14'd13038:data <=32'hFFE9FFCF;14'd13039:data <=32'hFFE3FFCF;14'd13040:data <=32'hFFDDFFCF;
14'd13041:data <=32'hFFD5FFD0;14'd13042:data <=32'hFFCBFFD3;14'd13043:data <=32'hFFC1FFD9;
14'd13044:data <=32'hFFB8FFE3;14'd13045:data <=32'hFFB3FFEF;14'd13046:data <=32'hFFB0FFFC;
14'd13047:data <=32'hFFB2000A;14'd13048:data <=32'hFFB60015;14'd13049:data <=32'hFFBC001F;
14'd13050:data <=32'hFFC30026;14'd13051:data <=32'hFFCA002C;14'd13052:data <=32'hFFD10030;
14'd13053:data <=32'hFFD90033;14'd13054:data <=32'hFFE10034;14'd13055:data <=32'hFFE80034;
14'd13056:data <=32'hFF9C003B;14'd13057:data <=32'hFFA30055;14'd13058:data <=32'hFFB90064;
14'd13059:data <=32'hFFEB0032;14'd13060:data <=32'hFFE80016;14'd13061:data <=32'hFFE00019;
14'd13062:data <=32'hFFDA0021;14'd13063:data <=32'hFFD6002D;14'd13064:data <=32'hFFD8003C;
14'd13065:data <=32'hFFE0004A;14'd13066:data <=32'hFFED0056;14'd13067:data <=32'hFFFE005D;
14'd13068:data <=32'h00100060;14'd13069:data <=32'h0022005E;14'd13070:data <=32'h00340057;
14'd13071:data <=32'h0043004E;14'd13072:data <=32'h00500040;14'd13073:data <=32'h005B0030;
14'd13074:data <=32'h0062001D;14'd13075:data <=32'h00640009;14'd13076:data <=32'h0061FFF5;
14'd13077:data <=32'h0058FFE2;14'd13078:data <=32'h004AFFD4;14'd13079:data <=32'h003AFFCA;
14'd13080:data <=32'h0028FFC6;14'd13081:data <=32'h0018FFC8;14'd13082:data <=32'h000BFFCD;
14'd13083:data <=32'h0002FFD5;14'd13084:data <=32'hFFFCFFDD;14'd13085:data <=32'hFFF9FFE4;
14'd13086:data <=32'hFFF8FFEB;14'd13087:data <=32'hFFF8FFF1;14'd13088:data <=32'hFFF8FFF7;
14'd13089:data <=32'hFFFAFFFE;14'd13090:data <=32'hFFFC0003;14'd13091:data <=32'h00020008;
14'd13092:data <=32'h0009000C;14'd13093:data <=32'h0011000D;14'd13094:data <=32'h001A000C;
14'd13095:data <=32'h00220007;14'd13096:data <=32'h00290001;14'd13097:data <=32'h002EFFF9;
14'd13098:data <=32'h0032FFEF;14'd13099:data <=32'h0034FFE5;14'd13100:data <=32'h0034FFDA;
14'd13101:data <=32'h0032FFCE;14'd13102:data <=32'h002DFFC1;14'd13103:data <=32'h0026FFB3;
14'd13104:data <=32'h0019FFA7;14'd13105:data <=32'h0008FF9D;14'd13106:data <=32'hFFF4FF97;
14'd13107:data <=32'hFFDEFF98;14'd13108:data <=32'hFFC7FF9F;14'd13109:data <=32'hFFB4FFAC;
14'd13110:data <=32'hFFA5FFBE;14'd13111:data <=32'hFF9CFFD2;14'd13112:data <=32'hFF99FFE7;
14'd13113:data <=32'hFF9BFFFA;14'd13114:data <=32'hFFA1000C;14'd13115:data <=32'hFFAB0019;
14'd13116:data <=32'hFFB50024;14'd13117:data <=32'hFFC1002B;14'd13118:data <=32'hFFCE002F;
14'd13119:data <=32'hFFDA0030;14'd13120:data <=32'hFFB8FFFE;14'd13121:data <=32'hFFB1000A;
14'd13122:data <=32'hFFB3001E;14'd13123:data <=32'hFFD90035;14'd13124:data <=32'hFFDE0017;
14'd13125:data <=32'hFFDB0015;14'd13126:data <=32'hFFD60017;14'd13127:data <=32'hFFD2001C;
14'd13128:data <=32'hFFD00025;14'd13129:data <=32'hFFD2002F;14'd13130:data <=32'hFFD80039;
14'd13131:data <=32'hFFE10041;14'd13132:data <=32'hFFEB0045;14'd13133:data <=32'hFFF60048;
14'd13134:data <=32'h00010048;14'd13135:data <=32'h000A0047;14'd13136:data <=32'h00140044;
14'd13137:data <=32'h001D0040;14'd13138:data <=32'h0025003A;14'd13139:data <=32'h002D0032;
14'd13140:data <=32'h00320029;14'd13141:data <=32'h0034001E;14'd13142:data <=32'h00350015;
14'd13143:data <=32'h0032000D;14'd13144:data <=32'h002E0006;14'd13145:data <=32'h002A0003;
14'd13146:data <=32'h00270001;14'd13147:data <=32'h0026FFFF;14'd13148:data <=32'h0025FFFC;
14'd13149:data <=32'h0024FFF9;14'd13150:data <=32'h0022FFF4;14'd13151:data <=32'h001FFFEF;
14'd13152:data <=32'h0019FFEB;14'd13153:data <=32'h0011FFEA;14'd13154:data <=32'h0009FFEB;
14'd13155:data <=32'h0003FFF0;14'd13156:data <=32'hFFFEFFF7;14'd13157:data <=32'hFFFCFFFF;
14'd13158:data <=32'hFFFE0008;14'd13159:data <=32'h0002000F;14'd13160:data <=32'h00090015;
14'd13161:data <=32'h00120019;14'd13162:data <=32'h001C001B;14'd13163:data <=32'h0028001A;
14'd13164:data <=32'h00340015;14'd13165:data <=32'h0040000D;14'd13166:data <=32'h004B0001;
14'd13167:data <=32'h0052FFF0;14'd13168:data <=32'h0055FFDC;14'd13169:data <=32'h0052FFC7;
14'd13170:data <=32'h0048FFB2;14'd13171:data <=32'h0038FFA1;14'd13172:data <=32'h0024FF95;
14'd13173:data <=32'h000EFF8F;14'd13174:data <=32'hFFF7FF8F;14'd13175:data <=32'hFFE3FF95;
14'd13176:data <=32'hFFD2FF9F;14'd13177:data <=32'hFFC5FFAB;14'd13178:data <=32'hFFBBFFB7;
14'd13179:data <=32'hFFB4FFC5;14'd13180:data <=32'hFFAFFFD1;14'd13181:data <=32'hFFADFFDF;
14'd13182:data <=32'hFFADFFEB;14'd13183:data <=32'hFFAFFFF6;14'd13184:data <=32'hFFC50000;
14'd13185:data <=32'hFFC60004;14'd13186:data <=32'hFFC10006;14'd13187:data <=32'hFFA40002;
14'd13188:data <=32'hFFA7FFF2;14'd13189:data <=32'hFFA4FFFD;14'd13190:data <=32'hFFA2000A;
14'd13191:data <=32'hFFA20019;14'd13192:data <=32'hFFA70029;14'd13193:data <=32'hFFAF0038;
14'd13194:data <=32'hFFBD0045;14'd13195:data <=32'hFFCD004E;14'd13196:data <=32'hFFDF0051;
14'd13197:data <=32'hFFF0004F;14'd13198:data <=32'hFFFE0049;14'd13199:data <=32'h00080041;
14'd13200:data <=32'h00100038;14'd13201:data <=32'h0014002F;14'd13202:data <=32'h00160026;
14'd13203:data <=32'h0016001F;14'd13204:data <=32'h00150018;14'd13205:data <=32'h00110012;
14'd13206:data <=32'h000C000F;14'd13207:data <=32'h0007000E;14'd13208:data <=32'h00010010;
14'd13209:data <=32'hFFFE0014;14'd13210:data <=32'hFFFE001B;14'd13211:data <=32'h00010021;
14'd13212:data <=32'h00070025;14'd13213:data <=32'h00100027;14'd13214:data <=32'h00180025;
14'd13215:data <=32'h0020001F;14'd13216:data <=32'h00240017;14'd13217:data <=32'h0024000F;
14'd13218:data <=32'h00220007;14'd13219:data <=32'h001E0002;14'd13220:data <=32'h00180000;
14'd13221:data <=32'h0014FFFF;14'd13222:data <=32'h000F0001;14'd13223:data <=32'h000C0004;
14'd13224:data <=32'h000B0007;14'd13225:data <=32'h000B000C;14'd13226:data <=32'h000C0010;
14'd13227:data <=32'h00100015;14'd13228:data <=32'h00160019;14'd13229:data <=32'h001D001B;
14'd13230:data <=32'h0027001C;14'd13231:data <=32'h00310018;14'd13232:data <=32'h003B0011;
14'd13233:data <=32'h00430007;14'd13234:data <=32'h0048FFFA;14'd13235:data <=32'h0048FFED;
14'd13236:data <=32'h0045FFE0;14'd13237:data <=32'h0040FFD5;14'd13238:data <=32'h0039FFCE;
14'd13239:data <=32'h0033FFC7;14'd13240:data <=32'h002CFFC2;14'd13241:data <=32'h0027FFBD;
14'd13242:data <=32'h0021FFB7;14'd13243:data <=32'h001AFFB0;14'd13244:data <=32'h0011FFA9;
14'd13245:data <=32'h0006FFA4;14'd13246:data <=32'hFFF9FFA0;14'd13247:data <=32'hFFEAFF9F;
14'd13248:data <=32'hFFC0FFD4;14'd13249:data <=32'hFFBFFFDC;14'd13250:data <=32'hFFC4FFDB;
14'd13251:data <=32'hFFD1FFA3;14'd13252:data <=32'hFFC2FF8E;14'd13253:data <=32'hFFABFF98;
14'd13254:data <=32'hFF97FFA9;14'd13255:data <=32'hFF86FFBE;14'd13256:data <=32'hFF7BFFD8;
14'd13257:data <=32'hFF77FFF6;14'd13258:data <=32'hFF7C0013;14'd13259:data <=32'hFF89002C;
14'd13260:data <=32'hFF9C0040;14'd13261:data <=32'hFFB1004D;14'd13262:data <=32'hFFC80053;
14'd13263:data <=32'hFFDC0053;14'd13264:data <=32'hFFEE004F;14'd13265:data <=32'hFFFD0047;
14'd13266:data <=32'h0009003D;14'd13267:data <=32'h00110032;14'd13268:data <=32'h00150026;
14'd13269:data <=32'h0016001A;14'd13270:data <=32'h0014000F;14'd13271:data <=32'h000D0006;
14'd13272:data <=32'h00050001;14'd13273:data <=32'hFFFC0000;14'd13274:data <=32'hFFF40003;
14'd13275:data <=32'hFFEE0009;14'd13276:data <=32'hFFED0010;14'd13277:data <=32'hFFEE0017;
14'd13278:data <=32'hFFF1001C;14'd13279:data <=32'hFFF5001F;14'd13280:data <=32'hFFFA0020;
14'd13281:data <=32'hFFFD0020;14'd13282:data <=32'hFFFF0020;14'd13283:data <=32'h00010020;
14'd13284:data <=32'h00020021;14'd13285:data <=32'h00040023;14'd13286:data <=32'h00080025;
14'd13287:data <=32'h000B0026;14'd13288:data <=32'h00110026;14'd13289:data <=32'h00160025;
14'd13290:data <=32'h001B0023;14'd13291:data <=32'h001E001F;14'd13292:data <=32'h0021001D;
14'd13293:data <=32'h0024001A;14'd13294:data <=32'h00270016;14'd13295:data <=32'h00290013;
14'd13296:data <=32'h002B000E;14'd13297:data <=32'h002C0009;14'd13298:data <=32'h002B0004;
14'd13299:data <=32'h002A0000;14'd13300:data <=32'h0026FFFD;14'd13301:data <=32'h0023FFFD;
14'd13302:data <=32'h0021FFFF;14'd13303:data <=32'h00220003;14'd13304:data <=32'h00270006;
14'd13305:data <=32'h002F0008;14'd13306:data <=32'h003A0005;14'd13307:data <=32'h0045FFFD;
14'd13308:data <=32'h004EFFF0;14'd13309:data <=32'h0053FFE0;14'd13310:data <=32'h0053FFCD;
14'd13311:data <=32'h004FFFBA;14'd13312:data <=32'h000EFFB5;14'd13313:data <=32'h0009FFB0;
14'd13314:data <=32'h000AFFB2;14'd13315:data <=32'h0034FFB0;14'd13316:data <=32'h002AFF88;
14'd13317:data <=32'h0013FF7E;14'd13318:data <=32'hFFF8FF7A;14'd13319:data <=32'hFFDEFF7D;
14'd13320:data <=32'hFFC4FF88;14'd13321:data <=32'hFFAEFF99;14'd13322:data <=32'hFF9EFFAF;
14'd13323:data <=32'hFF95FFC7;14'd13324:data <=32'hFF94FFDE;14'd13325:data <=32'hFF98FFF3;
14'd13326:data <=32'hFF9F0004;14'd13327:data <=32'hFFA90012;14'd13328:data <=32'hFFB3001C;
14'd13329:data <=32'hFFBD0024;14'd13330:data <=32'hFFC80029;14'd13331:data <=32'hFFD3002D;
14'd13332:data <=32'hFFDE002E;14'd13333:data <=32'hFFE8002D;14'd13334:data <=32'hFFF10029;
14'd13335:data <=32'hFFF80024;14'd13336:data <=32'hFFFC001E;14'd13337:data <=32'hFFFE0018;
14'd13338:data <=32'hFFFE0014;14'd13339:data <=32'hFFFE0011;14'd13340:data <=32'hFFFE000E;
14'd13341:data <=32'hFFFD000C;14'd13342:data <=32'hFFFD0009;14'd13343:data <=32'hFFFC0005;
14'd13344:data <=32'hFFF90001;14'd13345:data <=32'hFFF4FFFF;14'd13346:data <=32'hFFEDFFFE;
14'd13347:data <=32'hFFE50000;14'd13348:data <=32'hFFDE0005;14'd13349:data <=32'hFFD8000F;
14'd13350:data <=32'hFFD6001A;14'd13351:data <=32'hFFD80026;14'd13352:data <=32'hFFDD0031;
14'd13353:data <=32'hFFE6003A;14'd13354:data <=32'hFFF10040;14'd13355:data <=32'hFFFD0043;
14'd13356:data <=32'h00080043;14'd13357:data <=32'h00140042;14'd13358:data <=32'h001E003D;
14'd13359:data <=32'h00270036;14'd13360:data <=32'h002E002E;14'd13361:data <=32'h00340024;
14'd13362:data <=32'h00350019;14'd13363:data <=32'h0032000F;14'd13364:data <=32'h002E0007;
14'd13365:data <=32'h00260002;14'd13366:data <=32'h001F0002;14'd13367:data <=32'h00190006;
14'd13368:data <=32'h0017000C;14'd13369:data <=32'h001A0014;14'd13370:data <=32'h0021001A;
14'd13371:data <=32'h002B001D;14'd13372:data <=32'h0038001A;14'd13373:data <=32'h00440014;
14'd13374:data <=32'h004E0009;14'd13375:data <=32'h0055FFFC;14'd13376:data <=32'h00460002;
14'd13377:data <=32'h0054FFF5;14'd13378:data <=32'h0056FFEB;14'd13379:data <=32'h0042FFEC;
14'd13380:data <=32'h0045FFC6;14'd13381:data <=32'h003CFFBB;14'd13382:data <=32'h0030FFB2;
14'd13383:data <=32'h0022FFAB;14'd13384:data <=32'h0013FFA9;14'd13385:data <=32'h0004FFAA;
14'd13386:data <=32'hFFF8FFAF;14'd13387:data <=32'hFFEEFFB6;14'd13388:data <=32'hFFE8FFBD;
14'd13389:data <=32'hFFE4FFC3;14'd13390:data <=32'hFFE1FFC7;14'd13391:data <=32'hFFDEFFCA;
14'd13392:data <=32'hFFD9FFCC;14'd13393:data <=32'hFFD3FFCF;14'd13394:data <=32'hFFCCFFD4;
14'd13395:data <=32'hFFC6FFDC;14'd13396:data <=32'hFFC1FFE6;14'd13397:data <=32'hFFBFFFF0;
14'd13398:data <=32'hFFC0FFFA;14'd13399:data <=32'hFFC20004;14'd13400:data <=32'hFFC6000D;
14'd13401:data <=32'hFFCC0015;14'd13402:data <=32'hFFD2001C;14'd13403:data <=32'hFFDB0021;
14'd13404:data <=32'hFFE50025;14'd13405:data <=32'hFFF00025;14'd13406:data <=32'hFFFB0022;
14'd13407:data <=32'h0004001B;14'd13408:data <=32'h000B0011;14'd13409:data <=32'h000D0004;
14'd13410:data <=32'h000AFFF9;14'd13411:data <=32'h0002FFEE;14'd13412:data <=32'hFFF7FFE8;
14'd13413:data <=32'hFFEAFFE7;14'd13414:data <=32'hFFDDFFEA;14'd13415:data <=32'hFFD3FFF1;
14'd13416:data <=32'hFFCBFFFC;14'd13417:data <=32'hFFC70007;14'd13418:data <=32'hFFC50013;
14'd13419:data <=32'hFFC8001F;14'd13420:data <=32'hFFCB002A;14'd13421:data <=32'hFFD20034;
14'd13422:data <=32'hFFDA003C;14'd13423:data <=32'hFFE40043;14'd13424:data <=32'hFFEE0047;
14'd13425:data <=32'hFFFA0049;14'd13426:data <=32'h00050047;14'd13427:data <=32'h000F0043;
14'd13428:data <=32'h0016003F;14'd13429:data <=32'h001A003A;14'd13430:data <=32'h001D0036;
14'd13431:data <=32'h00200034;14'd13432:data <=32'h00230033;14'd13433:data <=32'h00280034;
14'd13434:data <=32'h00300033;14'd13435:data <=32'h00390030;14'd13436:data <=32'h0043002A;
14'd13437:data <=32'h004C0020;14'd13438:data <=32'h00520014;14'd13439:data <=32'h00540007;
14'd13440:data <=32'h0017003A;14'd13441:data <=32'h002E0040;14'd13442:data <=32'h00440036;
14'd13443:data <=32'h0045FFF3;14'd13444:data <=32'h0045FFD2;14'd13445:data <=32'h0039FFCC;
14'd13446:data <=32'h002CFFC8;14'd13447:data <=32'h0021FFC8;14'd13448:data <=32'h0016FFCA;
14'd13449:data <=32'h000DFFCF;14'd13450:data <=32'h0007FFD7;14'd13451:data <=32'h0006FFE0;
14'd13452:data <=32'h0009FFE6;14'd13453:data <=32'h000FFFE9;14'd13454:data <=32'h0015FFE8;
14'd13455:data <=32'h001AFFE2;14'd13456:data <=32'h001CFFD9;14'd13457:data <=32'h001AFFCF;
14'd13458:data <=32'h0013FFC5;14'd13459:data <=32'h0009FFBF;14'd13460:data <=32'hFFFDFFBB;
14'd13461:data <=32'hFFF0FFBB;14'd13462:data <=32'hFFE4FFBF;14'd13463:data <=32'hFFDAFFC5;
14'd13464:data <=32'hFFD1FFCD;14'd13465:data <=32'hFFC9FFD7;14'd13466:data <=32'hFFC4FFE3;
14'd13467:data <=32'hFFC2FFEF;14'd13468:data <=32'hFFC3FFFD;14'd13469:data <=32'hFFCA0009;
14'd13470:data <=32'hFFD30013;14'd13471:data <=32'hFFDE0019;14'd13472:data <=32'hFFEB001A;
14'd13473:data <=32'hFFF60016;14'd13474:data <=32'hFFFE000F;14'd13475:data <=32'h00030007;
14'd13476:data <=32'h0003FFFE;14'd13477:data <=32'h0001FFF6;14'd13478:data <=32'hFFFCFFF1;
14'd13479:data <=32'hFFF6FFED;14'd13480:data <=32'hFFF1FFEB;14'd13481:data <=32'hFFEBFFEA;
14'd13482:data <=32'hFFE5FFEB;14'd13483:data <=32'hFFDFFFEB;14'd13484:data <=32'hFFD9FFED;
14'd13485:data <=32'hFFD2FFF0;14'd13486:data <=32'hFFCAFFF5;14'd13487:data <=32'hFFC4FFFC;
14'd13488:data <=32'hFFBE0006;14'd13489:data <=32'hFFBB0010;14'd13490:data <=32'hFFBA001C;
14'd13491:data <=32'hFFBB0028;14'd13492:data <=32'hFFBE0034;14'd13493:data <=32'hFFC20040;
14'd13494:data <=32'hFFC9004C;14'd13495:data <=32'hFFD20059;14'd13496:data <=32'hFFDF0065;
14'd13497:data <=32'hFFF00070;14'd13498:data <=32'h00040077;14'd13499:data <=32'h001B0079;
14'd13500:data <=32'h00340074;14'd13501:data <=32'h004B0068;14'd13502:data <=32'h005E0056;
14'd13503:data <=32'h006B0040;14'd13504:data <=32'h0000002D;14'd13505:data <=32'h000B003C;
14'd13506:data <=32'h00230046;14'd13507:data <=32'h0065002A;14'd13508:data <=32'h006BFFFD;
14'd13509:data <=32'h0061FFEC;14'd13510:data <=32'h0054FFDE;14'd13511:data <=32'h0046FFD4;
14'd13512:data <=32'h0036FFCF;14'd13513:data <=32'h0027FFCF;14'd13514:data <=32'h001AFFD4;
14'd13515:data <=32'h0010FFDB;14'd13516:data <=32'h000DFFE5;14'd13517:data <=32'h000DFFED;
14'd13518:data <=32'h0012FFF3;14'd13519:data <=32'h0019FFF4;14'd13520:data <=32'h001FFFF2;
14'd13521:data <=32'h0023FFEC;14'd13522:data <=32'h0023FFE5;14'd13523:data <=32'h0021FFDE;
14'd13524:data <=32'h001DFFD7;14'd13525:data <=32'h0017FFD3;14'd13526:data <=32'h0011FFD0;
14'd13527:data <=32'h000BFFCE;14'd13528:data <=32'h0004FFCD;14'd13529:data <=32'hFFFEFFCD;
14'd13530:data <=32'hFFF7FFCF;14'd13531:data <=32'hFFF0FFD2;14'd13532:data <=32'hFFE9FFD7;
14'd13533:data <=32'hFFE5FFDD;14'd13534:data <=32'hFFE3FFE4;14'd13535:data <=32'hFFE4FFEA;
14'd13536:data <=32'hFFE6FFEF;14'd13537:data <=32'hFFE9FFF2;14'd13538:data <=32'hFFEBFFF4;
14'd13539:data <=32'hFFECFFF4;14'd13540:data <=32'hFFEDFFF4;14'd13541:data <=32'hFFECFFF5;
14'd13542:data <=32'hFFECFFF7;14'd13543:data <=32'hFFEDFFF9;14'd13544:data <=32'hFFF0FFFC;
14'd13545:data <=32'hFFF3FFFC;14'd13546:data <=32'hFFF8FFFB;14'd13547:data <=32'hFFFCFFF7;
14'd13548:data <=32'hFFFFFFF0;14'd13549:data <=32'hFFFEFFE8;14'd13550:data <=32'hFFFAFFDF;
14'd13551:data <=32'hFFF2FFD8;14'd13552:data <=32'hFFE7FFD3;14'd13553:data <=32'hFFDAFFD1;
14'd13554:data <=32'hFFCCFFD2;14'd13555:data <=32'hFFBEFFD8;14'd13556:data <=32'hFFB0FFE0;
14'd13557:data <=32'hFFA3FFED;14'd13558:data <=32'hFF98FFFD;14'd13559:data <=32'hFF910012;
14'd13560:data <=32'hFF8E002A;14'd13561:data <=32'hFF920044;14'd13562:data <=32'hFF9E005D;
14'd13563:data <=32'hFFB10074;14'd13564:data <=32'hFFCA0084;14'd13565:data <=32'hFFE7008D;
14'd13566:data <=32'h0005008E;14'd13567:data <=32'h00200087;14'd13568:data <=32'hFFFD004C;
14'd13569:data <=32'h00080056;14'd13570:data <=32'h00110063;14'd13571:data <=32'h00240079;
14'd13572:data <=32'h003C0055;14'd13573:data <=32'h00450048;14'd13574:data <=32'h004B003A;
14'd13575:data <=32'h004E002D;14'd13576:data <=32'h004F001F;14'd13577:data <=32'h004C0013;
14'd13578:data <=32'h0048000A;14'd13579:data <=32'h00440003;14'd13580:data <=32'h003FFFFF;
14'd13581:data <=32'h003DFFFB;14'd13582:data <=32'h003CFFF6;14'd13583:data <=32'h003BFFF1;
14'd13584:data <=32'h003AFFE9;14'd13585:data <=32'h0036FFE1;14'd13586:data <=32'h002FFFDA;
14'd13587:data <=32'h0026FFD5;14'd13588:data <=32'h001CFFD2;14'd13589:data <=32'h0012FFD4;
14'd13590:data <=32'h000AFFD8;14'd13591:data <=32'h0004FFDD;14'd13592:data <=32'h0002FFE3;
14'd13593:data <=32'h0001FFE8;14'd13594:data <=32'h0001FFEC;14'd13595:data <=32'h0003FFEF;
14'd13596:data <=32'h0005FFF1;14'd13597:data <=32'h0008FFF2;14'd13598:data <=32'h000AFFF2;
14'd13599:data <=32'h000DFFF1;14'd13600:data <=32'h0010FFED;14'd13601:data <=32'h0012FFE9;
14'd13602:data <=32'h0011FFE3;14'd13603:data <=32'h000EFFDD;14'd13604:data <=32'h0008FFD8;
14'd13605:data <=32'h0001FFD6;14'd13606:data <=32'hFFF8FFD6;14'd13607:data <=32'hFFF1FFDA;
14'd13608:data <=32'hFFECFFE0;14'd13609:data <=32'hFFEBFFE7;14'd13610:data <=32'hFFEDFFEE;
14'd13611:data <=32'hFFF1FFF2;14'd13612:data <=32'hFFF7FFF3;14'd13613:data <=32'hFFFCFFF1;
14'd13614:data <=32'h0000FFEC;14'd13615:data <=32'h0000FFE4;14'd13616:data <=32'hFFFFFFDD;
14'd13617:data <=32'hFFFAFFD6;14'd13618:data <=32'hFFF3FFD0;14'd13619:data <=32'hFFEAFFCB;
14'd13620:data <=32'hFFDFFFC9;14'd13621:data <=32'hFFD2FFC8;14'd13622:data <=32'hFFC4FFCB;
14'd13623:data <=32'hFFB5FFD2;14'd13624:data <=32'hFFA7FFDE;14'd13625:data <=32'hFF9CFFEE;
14'd13626:data <=32'hFF950002;14'd13627:data <=32'hFF950018;14'd13628:data <=32'hFF9A002D;
14'd13629:data <=32'hFFA5003E;14'd13630:data <=32'hFFB3004C;14'd13631:data <=32'hFFC20055;
14'd13632:data <=32'hFFB00057;14'd13633:data <=32'hFFBC006B;14'd13634:data <=32'hFFC70074;
14'd13635:data <=32'hFFC10053;14'd13636:data <=32'hFFD30043;14'd13637:data <=32'hFFD9004A;
14'd13638:data <=32'hFFE10051;14'd13639:data <=32'hFFEC0058;14'd13640:data <=32'hFFF8005C;
14'd13641:data <=32'h0006005F;14'd13642:data <=32'h0013005E;14'd13643:data <=32'h0021005D;
14'd13644:data <=32'h002F0059;14'd13645:data <=32'h003E0052;14'd13646:data <=32'h004D0047;
14'd13647:data <=32'h005A0039;14'd13648:data <=32'h00630026;14'd13649:data <=32'h00670010;
14'd13650:data <=32'h0064FFFA;14'd13651:data <=32'h005BFFE6;14'd13652:data <=32'h004DFFD6;
14'd13653:data <=32'h003CFFCC;14'd13654:data <=32'h002AFFC8;14'd13655:data <=32'h0019FFC9;
14'd13656:data <=32'h000BFFCE;14'd13657:data <=32'h0001FFD6;14'd13658:data <=32'hFFF9FFE0;
14'd13659:data <=32'hFFF5FFEA;14'd13660:data <=32'hFFF4FFF4;14'd13661:data <=32'hFFF6FFFD;
14'd13662:data <=32'hFFFB0005;14'd13663:data <=32'h0002000B;14'd13664:data <=32'h000B000F;
14'd13665:data <=32'h0015000E;14'd13666:data <=32'h001E000A;14'd13667:data <=32'h00250003;
14'd13668:data <=32'h0029FFFA;14'd13669:data <=32'h0029FFF1;14'd13670:data <=32'h0027FFE8;
14'd13671:data <=32'h0022FFE2;14'd13672:data <=32'h001DFFDE;14'd13673:data <=32'h0018FFDC;
14'd13674:data <=32'h0015FFDB;14'd13675:data <=32'h0013FFDA;14'd13676:data <=32'h0012FFD8;
14'd13677:data <=32'h0010FFD4;14'd13678:data <=32'h000DFFCF;14'd13679:data <=32'h0009FFCA;
14'd13680:data <=32'h0002FFC7;14'd13681:data <=32'hFFFAFFC4;14'd13682:data <=32'hFFF2FFC4;
14'd13683:data <=32'hFFE9FFC5;14'd13684:data <=32'hFFE2FFC7;14'd13685:data <=32'hFFDAFFCA;
14'd13686:data <=32'hFFD3FFCE;14'd13687:data <=32'hFFCCFFD3;14'd13688:data <=32'hFFC6FFDA;
14'd13689:data <=32'hFFC0FFE2;14'd13690:data <=32'hFFBDFFEC;14'd13691:data <=32'hFFBCFFF7;
14'd13692:data <=32'hFFBF0000;14'd13693:data <=32'hFFC30007;14'd13694:data <=32'hFFC9000C;
14'd13695:data <=32'hFFCD000D;14'd13696:data <=32'hFF8AFFFE;14'd13697:data <=32'hFF830015;
14'd13698:data <=32'hFF8B0029;14'd13699:data <=32'hFFC3000A;14'd13700:data <=32'hFFC8FFF6;
14'd13701:data <=32'hFFBDFFFD;14'd13702:data <=32'hFFB50008;14'd13703:data <=32'hFFB00016;
14'd13704:data <=32'hFFAF0025;14'd13705:data <=32'hFFB20035;14'd13706:data <=32'hFFB80046;
14'd13707:data <=32'hFFC30055;14'd13708:data <=32'hFFD10062;14'd13709:data <=32'hFFE3006D;
14'd13710:data <=32'hFFF90073;14'd13711:data <=32'h00110074;14'd13712:data <=32'h0029006D;
14'd13713:data <=32'h003E0060;14'd13714:data <=32'h004E004D;14'd13715:data <=32'h00570037;
14'd13716:data <=32'h005B0021;14'd13717:data <=32'h0057000D;14'd13718:data <=32'h004FFFFD;
14'd13719:data <=32'h0045FFF0;14'd13720:data <=32'h0038FFE8;14'd13721:data <=32'h002DFFE3;
14'd13722:data <=32'h0022FFE0;14'd13723:data <=32'h0017FFE0;14'd13724:data <=32'h000DFFE2;
14'd13725:data <=32'h0004FFE7;14'd13726:data <=32'hFFFEFFED;14'd13727:data <=32'hFFF9FFF6;
14'd13728:data <=32'hFFF8FFFF;14'd13729:data <=32'hFFFA0007;14'd13730:data <=32'hFFFE000F;
14'd13731:data <=32'h00040013;14'd13732:data <=32'h000B0016;14'd13733:data <=32'h00110017;
14'd13734:data <=32'h00180017;14'd13735:data <=32'h001E0016;14'd13736:data <=32'h00250015;
14'd13737:data <=32'h002C0012;14'd13738:data <=32'h0034000E;14'd13739:data <=32'h003D0008;
14'd13740:data <=32'h0044FFFE;14'd13741:data <=32'h004AFFF0;14'd13742:data <=32'h004CFFE0;
14'd13743:data <=32'h0049FFCE;14'd13744:data <=32'h0041FFBD;14'd13745:data <=32'h0035FFB0;
14'd13746:data <=32'h0025FFA5;14'd13747:data <=32'h0013FF9F;14'd13748:data <=32'h0001FF9E;
14'd13749:data <=32'hFFF0FFA0;14'd13750:data <=32'hFFE0FFA7;14'd13751:data <=32'hFFD2FFAF;
14'd13752:data <=32'hFFC7FFBB;14'd13753:data <=32'hFFBEFFC8;14'd13754:data <=32'hFFBAFFD7;
14'd13755:data <=32'hFFB9FFE7;14'd13756:data <=32'hFFBEFFF4;14'd13757:data <=32'hFFC6FFFF;
14'd13758:data <=32'hFFD10005;14'd13759:data <=32'hFFDB0005;14'd13760:data <=32'hFFCAFFCC;
14'd13761:data <=32'hFFBCFFCE;14'd13762:data <=32'hFFB2FFDE;14'd13763:data <=32'hFFCE0000;
14'd13764:data <=32'hFFD8FFE7;14'd13765:data <=32'hFFD1FFE7;14'd13766:data <=32'hFFC8FFEA;
14'd13767:data <=32'hFFC0FFF1;14'd13768:data <=32'hFFBBFFFA;14'd13769:data <=32'hFFB70003;
14'd13770:data <=32'hFFB5000E;14'd13771:data <=32'hFFB5001A;14'd13772:data <=32'hFFB70027;
14'd13773:data <=32'hFFBC0034;14'd13774:data <=32'hFFC50040;14'd13775:data <=32'hFFD2004A;
14'd13776:data <=32'hFFE10050;14'd13777:data <=32'hFFF10052;14'd13778:data <=32'h0000004F;
14'd13779:data <=32'h000C0048;14'd13780:data <=32'h00150040;14'd13781:data <=32'h001B0037;
14'd13782:data <=32'h001E0030;14'd13783:data <=32'h0020002A;14'd13784:data <=32'h00210024;
14'd13785:data <=32'h00230020;14'd13786:data <=32'h0025001A;14'd13787:data <=32'h00270014;
14'd13788:data <=32'h0027000D;14'd13789:data <=32'h00250006;14'd13790:data <=32'h00210000;
14'd13791:data <=32'h001BFFFB;14'd13792:data <=32'h0015FFF8;14'd13793:data <=32'h000EFFF8;
14'd13794:data <=32'h0009FFF9;14'd13795:data <=32'h0003FFFB;14'd13796:data <=32'hFFFFFFFF;
14'd13797:data <=32'hFFFB0004;14'd13798:data <=32'hFFF8000B;14'd13799:data <=32'hFFF70014;
14'd13800:data <=32'hFFF9001E;14'd13801:data <=32'hFFFE0028;14'd13802:data <=32'h00080032;
14'd13803:data <=32'h00170038;14'd13804:data <=32'h0028003A;14'd13805:data <=32'h003A0036;
14'd13806:data <=32'h004C002C;14'd13807:data <=32'h005A001C;14'd13808:data <=32'h00630009;
14'd13809:data <=32'h0066FFF3;14'd13810:data <=32'h0064FFDE;14'd13811:data <=32'h005CFFCB;
14'd13812:data <=32'h0051FFBB;14'd13813:data <=32'h0043FFAD;14'd13814:data <=32'h0033FFA4;
14'd13815:data <=32'h0022FF9E;14'd13816:data <=32'h0010FF9B;14'd13817:data <=32'hFFFFFF9D;
14'd13818:data <=32'hFFEFFFA3;14'd13819:data <=32'hFFE1FFAC;14'd13820:data <=32'hFFD8FFB8;
14'd13821:data <=32'hFFD3FFC4;14'd13822:data <=32'hFFD2FFCF;14'd13823:data <=32'hFFD4FFD6;
14'd13824:data <=32'hFFE6FFE3;14'd13825:data <=32'hFFE7FFDE;14'd13826:data <=32'hFFDFFFD9;
14'd13827:data <=32'hFFC1FFCE;14'd13828:data <=32'hFFC6FFBE;14'd13829:data <=32'hFFBCFFC6;
14'd13830:data <=32'hFFB3FFD2;14'd13831:data <=32'hFFACFFE0;14'd13832:data <=32'hFFAAFFEF;
14'd13833:data <=32'hFFACFFFD;14'd13834:data <=32'hFFB0000A;14'd13835:data <=32'hFFB60014;
14'd13836:data <=32'hFFBD001D;14'd13837:data <=32'hFFC50024;14'd13838:data <=32'hFFCE002A;
14'd13839:data <=32'hFFD8002D;14'd13840:data <=32'hFFE3002E;14'd13841:data <=32'hFFEC002C;
14'd13842:data <=32'hFFF40027;14'd13843:data <=32'hFFF80020;14'd13844:data <=32'hFFF90019;
14'd13845:data <=32'hFFF70014;14'd13846:data <=32'hFFF20012;14'd13847:data <=32'hFFEE0013;
14'd13848:data <=32'hFFEA0018;14'd13849:data <=32'hFFEA001E;14'd13850:data <=32'hFFED0025;
14'd13851:data <=32'hFFF3002A;14'd13852:data <=32'hFFFA002C;14'd13853:data <=32'h0002002C;
14'd13854:data <=32'h0009002A;14'd13855:data <=32'h000F0026;14'd13856:data <=32'h00130020;
14'd13857:data <=32'h0015001B;14'd13858:data <=32'h00170015;14'd13859:data <=32'h0015000F;
14'd13860:data <=32'h00130009;14'd13861:data <=32'h000F0005;14'd13862:data <=32'h00080003;
14'd13863:data <=32'h00010003;14'd13864:data <=32'hFFFA0007;14'd13865:data <=32'hFFF4000F;
14'd13866:data <=32'hFFF20019;14'd13867:data <=32'hFFF40024;14'd13868:data <=32'hFFFB002E;
14'd13869:data <=32'h00050036;14'd13870:data <=32'h0012003B;14'd13871:data <=32'h0020003A;
14'd13872:data <=32'h002D0037;14'd13873:data <=32'h0039002F;14'd13874:data <=32'h00410026;
14'd13875:data <=32'h0047001D;14'd13876:data <=32'h004C0013;14'd13877:data <=32'h004F0009;
14'd13878:data <=32'h0052FFFE;14'd13879:data <=32'h0052FFF3;14'd13880:data <=32'h0052FFE7;
14'd13881:data <=32'h0050FFDB;14'd13882:data <=32'h004BFFD0;14'd13883:data <=32'h0045FFC6;
14'd13884:data <=32'h003DFFBD;14'd13885:data <=32'h0035FFB6;14'd13886:data <=32'h002DFFAF;
14'd13887:data <=32'h0025FFA8;14'd13888:data <=32'hFFEBFFCF;14'd13889:data <=32'hFFEEFFD2;
14'd13890:data <=32'hFFF5FFCC;14'd13891:data <=32'h000FFF94;14'd13892:data <=32'h0007FF79;
14'd13893:data <=32'hFFEBFF79;14'd13894:data <=32'hFFD0FF80;14'd13895:data <=32'hFFB8FF8F;
14'd13896:data <=32'hFFA6FFA3;14'd13897:data <=32'hFF9AFFBA;14'd13898:data <=32'hFF95FFD2;
14'd13899:data <=32'hFF95FFE8;14'd13900:data <=32'hFF9AFFFD;14'd13901:data <=32'hFFA2000F;
14'd13902:data <=32'hFFAF001E;14'd13903:data <=32'hFFBD0029;14'd13904:data <=32'hFFCD002F;
14'd13905:data <=32'hFFDE0031;14'd13906:data <=32'hFFED002D;14'd13907:data <=32'hFFF90024;
14'd13908:data <=32'h00000019;14'd13909:data <=32'h0002000E;14'd13910:data <=32'hFFFF0004;
14'd13911:data <=32'hFFF8FFFD;14'd13912:data <=32'hFFF1FFFB;14'd13913:data <=32'hFFE9FFFC;
14'd13914:data <=32'hFFE40001;14'd13915:data <=32'hFFE10006;14'd13916:data <=32'hFFE1000C;
14'd13917:data <=32'hFFE20011;14'd13918:data <=32'hFFE40015;14'd13919:data <=32'hFFE60017;
14'd13920:data <=32'hFFE8001A;14'd13921:data <=32'hFFEB001D;14'd13922:data <=32'hFFEE001F;
14'd13923:data <=32'hFFF10020;14'd13924:data <=32'hFFF50021;14'd13925:data <=32'hFFF80020;
14'd13926:data <=32'hFFFB001F;14'd13927:data <=32'hFFFC001E;14'd13928:data <=32'hFFFC001D;
14'd13929:data <=32'hFFFC001D;14'd13930:data <=32'hFFFC001F;14'd13931:data <=32'hFFFD0022;
14'd13932:data <=32'h00000025;14'd13933:data <=32'h00040028;14'd13934:data <=32'h00090028;
14'd13935:data <=32'h000E0026;14'd13936:data <=32'h00120024;14'd13937:data <=32'h00130021;
14'd13938:data <=32'h0014001E;14'd13939:data <=32'h0012001E;14'd13940:data <=32'h00110020;
14'd13941:data <=32'h00120024;14'd13942:data <=32'h00160029;14'd13943:data <=32'h001C002E;
14'd13944:data <=32'h00260031;14'd13945:data <=32'h00310031;14'd13946:data <=32'h003E002F;
14'd13947:data <=32'h004A0029;14'd13948:data <=32'h00570020;14'd13949:data <=32'h00620014;
14'd13950:data <=32'h006B0005;14'd13951:data <=32'h0073FFF2;14'd13952:data <=32'h002FFFD4;
14'd13953:data <=32'h0032FFCF;14'd13954:data <=32'h0039FFCF;14'd13955:data <=32'h0069FFD3;
14'd13956:data <=32'h006DFFA5;14'd13957:data <=32'h0058FF90;14'd13958:data <=32'h003EFF82;
14'd13959:data <=32'h0022FF7A;14'd13960:data <=32'h0007FF7B;14'd13961:data <=32'hFFEFFF82;
14'd13962:data <=32'hFFDAFF8E;14'd13963:data <=32'hFFCAFF9C;14'd13964:data <=32'hFFBDFFAC;
14'd13965:data <=32'hFFB5FFBD;14'd13966:data <=32'hFFB0FFCF;14'd13967:data <=32'hFFAFFFE0;
14'd13968:data <=32'hFFB3FFF0;14'd13969:data <=32'hFFBAFFFF;14'd13970:data <=32'hFFC40009;
14'd13971:data <=32'hFFCF000F;14'd13972:data <=32'hFFD90011;14'd13973:data <=32'hFFE10010;
14'd13974:data <=32'hFFE6000D;14'd13975:data <=32'hFFE9000A;14'd13976:data <=32'hFFEB0009;
14'd13977:data <=32'hFFEC0008;14'd13978:data <=32'hFFEE0008;14'd13979:data <=32'hFFF10008;
14'd13980:data <=32'hFFF30007;14'd13981:data <=32'hFFF60004;14'd13982:data <=32'hFFF70000;
14'd13983:data <=32'hFFF6FFFA;14'd13984:data <=32'hFFF2FFF7;14'd13985:data <=32'hFFECFFF4;
14'd13986:data <=32'hFFE6FFF4;14'd13987:data <=32'hFFE0FFF7;14'd13988:data <=32'hFFDAFFFB;
14'd13989:data <=32'hFFD60001;14'd13990:data <=32'hFFD20007;14'd13991:data <=32'hFFD1000F;
14'd13992:data <=32'hFFD10017;14'd13993:data <=32'hFFD3001F;14'd13994:data <=32'hFFD60028;
14'd13995:data <=32'hFFDB0030;14'd13996:data <=32'hFFE40037;14'd13997:data <=32'hFFEE003B;
14'd13998:data <=32'hFFFA003C;14'd13999:data <=32'h00050039;14'd14000:data <=32'h000E0032;
14'd14001:data <=32'h0013002A;14'd14002:data <=32'h00140021;14'd14003:data <=32'h0011001A;
14'd14004:data <=32'h000B0015;14'd14005:data <=32'h00040016;14'd14006:data <=32'hFFFF001A;
14'd14007:data <=32'hFFFC0021;14'd14008:data <=32'hFFFD002A;14'd14009:data <=32'h00000033;
14'd14010:data <=32'h0008003B;14'd14011:data <=32'h00130041;14'd14012:data <=32'h001F0045;
14'd14013:data <=32'h002E0047;14'd14014:data <=32'h003E0045;14'd14015:data <=32'h0050003E;
14'd14016:data <=32'h003E0030;14'd14017:data <=32'h0053002D;14'd14018:data <=32'h005D0026;
14'd14019:data <=32'h00530023;14'd14020:data <=32'h0068FFFD;14'd14021:data <=32'h0064FFEA;
14'd14022:data <=32'h005DFFDA;14'd14023:data <=32'h0052FFCD;14'd14024:data <=32'h0046FFC4;
14'd14025:data <=32'h003AFFBF;14'd14026:data <=32'h0030FFBC;14'd14027:data <=32'h0027FFB9;
14'd14028:data <=32'h001EFFB7;14'd14029:data <=32'h0015FFB5;14'd14030:data <=32'h000CFFB4;
14'd14031:data <=32'h0002FFB5;14'd14032:data <=32'hFFF8FFB7;14'd14033:data <=32'hFFEFFFBB;
14'd14034:data <=32'hFFE8FFC0;14'd14035:data <=32'hFFE1FFC6;14'd14036:data <=32'hFFDCFFCB;
14'd14037:data <=32'hFFD7FFD1;14'd14038:data <=32'hFFD2FFD7;14'd14039:data <=32'hFFCDFFDF;
14'd14040:data <=32'hFFC9FFE9;14'd14041:data <=32'hFFC8FFF5;14'd14042:data <=32'hFFCB0001;
14'd14043:data <=32'hFFD2000C;14'd14044:data <=32'hFFDC0014;14'd14045:data <=32'hFFE90017;
14'd14046:data <=32'hFFF50016;14'd14047:data <=32'h00000010;14'd14048:data <=32'h00060007;
14'd14049:data <=32'h0009FFFD;14'd14050:data <=32'h0008FFF3;14'd14051:data <=32'h0004FFE9;
14'd14052:data <=32'hFFFCFFE2;14'd14053:data <=32'hFFF4FFDE;14'd14054:data <=32'hFFEAFFDC;
14'd14055:data <=32'hFFDFFFDC;14'd14056:data <=32'hFFD5FFDF;14'd14057:data <=32'hFFCBFFE6;
14'd14058:data <=32'hFFC3FFEF;14'd14059:data <=32'hFFBDFFFB;14'd14060:data <=32'hFFBB0009;
14'd14061:data <=32'hFFBD0016;14'd14062:data <=32'hFFC20022;14'd14063:data <=32'hFFCB002B;
14'd14064:data <=32'hFFD50030;14'd14065:data <=32'hFFDE0032;14'd14066:data <=32'hFFE50032;
14'd14067:data <=32'hFFEA0030;14'd14068:data <=32'hFFEC002F;14'd14069:data <=32'hFFED0030;
14'd14070:data <=32'hFFEE0032;14'd14071:data <=32'hFFF00036;14'd14072:data <=32'hFFF4003B;
14'd14073:data <=32'hFFFA0040;14'd14074:data <=32'h00020043;14'd14075:data <=32'h000B0045;
14'd14076:data <=32'h00130045;14'd14077:data <=32'h001C0045;14'd14078:data <=32'h00260043;
14'd14079:data <=32'h00300040;14'd14080:data <=32'hFFEE0053;14'd14081:data <=32'h00040066;
14'd14082:data <=32'h001F0068;14'd14083:data <=32'h0037002B;14'd14084:data <=32'h004A000C;
14'd14085:data <=32'h00440000;14'd14086:data <=32'h003CFFF8;14'd14087:data <=32'h0033FFF3;
14'd14088:data <=32'h002AFFF3;14'd14089:data <=32'h0025FFF6;14'd14090:data <=32'h0024FFFB;
14'd14091:data <=32'h0026FFFE;14'd14092:data <=32'h002BFFFF;14'd14093:data <=32'h0031FFFC;
14'd14094:data <=32'h0036FFF7;14'd14095:data <=32'h0039FFEF;14'd14096:data <=32'h003AFFE5;
14'd14097:data <=32'h0039FFDB;14'd14098:data <=32'h0035FFD2;14'd14099:data <=32'h0030FFC8;
14'd14100:data <=32'h0027FFBF;14'd14101:data <=32'h001CFFB7;14'd14102:data <=32'h000FFFB1;
14'd14103:data <=32'hFFFEFFB0;14'd14104:data <=32'hFFEEFFB3;14'd14105:data <=32'hFFDFFFBB;
14'd14106:data <=32'hFFD3FFC8;14'd14107:data <=32'hFFCCFFD7;14'd14108:data <=32'hFFCBFFE7;
14'd14109:data <=32'hFFCFFFF6;14'd14110:data <=32'hFFD70001;14'd14111:data <=32'hFFE10009;
14'd14112:data <=32'hFFEC000B;14'd14113:data <=32'hFFF5000B;14'd14114:data <=32'hFFFD0007;
14'd14115:data <=32'h00030003;14'd14116:data <=32'h0008FFFC;14'd14117:data <=32'h000AFFF6;
14'd14118:data <=32'h000BFFEE;14'd14119:data <=32'h0009FFE6;14'd14120:data <=32'h0005FFDF;
14'd14121:data <=32'hFFFFFFD8;14'd14122:data <=32'hFFF7FFD3;14'd14123:data <=32'hFFEDFFD1;
14'd14124:data <=32'hFFE3FFD1;14'd14125:data <=32'hFFD9FFD3;14'd14126:data <=32'hFFD1FFD8;
14'd14127:data <=32'hFFCAFFDD;14'd14128:data <=32'hFFC4FFE3;14'd14129:data <=32'hFFBEFFEA;
14'd14130:data <=32'hFFB8FFF0;14'd14131:data <=32'hFFB2FFF8;14'd14132:data <=32'hFFAB0003;
14'd14133:data <=32'hFFA60010;14'd14134:data <=32'hFFA40020;14'd14135:data <=32'hFFA60033;
14'd14136:data <=32'hFFAC0046;14'd14137:data <=32'hFFB90057;14'd14138:data <=32'hFFCA0064;
14'd14139:data <=32'hFFDD006C;14'd14140:data <=32'hFFF10070;14'd14141:data <=32'h00050070;
14'd14142:data <=32'h0018006B;14'd14143:data <=32'h00290063;14'd14144:data <=32'hFFCF002B;
14'd14145:data <=32'hFFD30044;14'd14146:data <=32'hFFE7005B;14'd14147:data <=32'h00350055;
14'd14148:data <=32'h004F0030;14'd14149:data <=32'h004D001C;14'd14150:data <=32'h0046000C;
14'd14151:data <=32'h003B0000;14'd14152:data <=32'h002EFFFA;14'd14153:data <=32'h0023FFFA;
14'd14154:data <=32'h001BFFFF;14'd14155:data <=32'h00170006;14'd14156:data <=32'h0017000C;
14'd14157:data <=32'h001B0010;14'd14158:data <=32'h00200012;14'd14159:data <=32'h00270012;
14'd14160:data <=32'h002D000F;14'd14161:data <=32'h0032000A;14'd14162:data <=32'h00370004;
14'd14163:data <=32'h003AFFFC;14'd14164:data <=32'h003CFFF3;14'd14165:data <=32'h003CFFE9;
14'd14166:data <=32'h0038FFDD;14'd14167:data <=32'h0032FFD3;14'd14168:data <=32'h0027FFCB;
14'd14169:data <=32'h001CFFC7;14'd14170:data <=32'h000FFFC6;14'd14171:data <=32'h0004FFCA;
14'd14172:data <=32'hFFFCFFD0;14'd14173:data <=32'hFFF7FFD6;14'd14174:data <=32'hFFF4FFDD;
14'd14175:data <=32'hFFF3FFE2;14'd14176:data <=32'hFFF4FFE6;14'd14177:data <=32'hFFF4FFE9;
14'd14178:data <=32'hFFF4FFEC;14'd14179:data <=32'hFFF4FFEF;14'd14180:data <=32'hFFF4FFF2;
14'd14181:data <=32'hFFF6FFF5;14'd14182:data <=32'hFFF9FFF9;14'd14183:data <=32'hFFFEFFFB;
14'd14184:data <=32'h0003FFFB;14'd14185:data <=32'h0009FFF8;14'd14186:data <=32'h000DFFF4;
14'd14187:data <=32'h0011FFEE;14'd14188:data <=32'h0012FFE6;14'd14189:data <=32'h0012FFDE;
14'd14190:data <=32'h0010FFD6;14'd14191:data <=32'h000CFFCD;14'd14192:data <=32'h0005FFC3;
14'd14193:data <=32'hFFFBFFBA;14'd14194:data <=32'hFFEEFFB2;14'd14195:data <=32'hFFDDFFAD;
14'd14196:data <=32'hFFC8FFAD;14'd14197:data <=32'hFFB2FFB2;14'd14198:data <=32'hFF9CFFBF;
14'd14199:data <=32'hFF8AFFD3;14'd14200:data <=32'hFF7EFFEC;14'd14201:data <=32'hFF790007;
14'd14202:data <=32'hFF7C0023;14'd14203:data <=32'hFF85003E;14'd14204:data <=32'hFF940053;
14'd14205:data <=32'hFFA80065;14'd14206:data <=32'hFFBD0072;14'd14207:data <=32'hFFD50079;
14'd14208:data <=32'hFFCD0030;14'd14209:data <=32'hFFCD0041;14'd14210:data <=32'hFFCF0056;
14'd14211:data <=32'hFFE0007A;14'd14212:data <=32'h00070063;14'd14213:data <=32'h00150059;
14'd14214:data <=32'h001E004D;14'd14215:data <=32'h00230042;14'd14216:data <=32'h00240039;
14'd14217:data <=32'h00240032;14'd14218:data <=32'h0025002F;14'd14219:data <=32'h0026002C;
14'd14220:data <=32'h0029002A;14'd14221:data <=32'h002E0026;14'd14222:data <=32'h00320020;
14'd14223:data <=32'h00350019;14'd14224:data <=32'h00360011;14'd14225:data <=32'h00350009;
14'd14226:data <=32'h00330003;14'd14227:data <=32'h0030FFFE;14'd14228:data <=32'h002DFFFA;
14'd14229:data <=32'h0029FFF6;14'd14230:data <=32'h0026FFF3;14'd14231:data <=32'h0022FFF0;
14'd14232:data <=32'h001EFFEE;14'd14233:data <=32'h0019FFEE;14'd14234:data <=32'h0014FFEF;
14'd14235:data <=32'h0012FFF2;14'd14236:data <=32'h0010FFF6;14'd14237:data <=32'h0012FFF8;
14'd14238:data <=32'h0016FFFA;14'd14239:data <=32'h001AFFF9;14'd14240:data <=32'h001DFFF5;
14'd14241:data <=32'h001FFFEE;14'd14242:data <=32'h001DFFE8;14'd14243:data <=32'h0019FFE2;
14'd14244:data <=32'h0013FFDF;14'd14245:data <=32'h000BFFDF;14'd14246:data <=32'h0006FFE1;
14'd14247:data <=32'h0001FFE5;14'd14248:data <=32'h0000FFEA;14'd14249:data <=32'h0000FFEF;
14'd14250:data <=32'h0003FFF3;14'd14251:data <=32'h0006FFF5;14'd14252:data <=32'h000BFFF6;
14'd14253:data <=32'h0010FFF5;14'd14254:data <=32'h0016FFF1;14'd14255:data <=32'h001BFFEC;
14'd14256:data <=32'h0020FFE4;14'd14257:data <=32'h0022FFD8;14'd14258:data <=32'h0021FFCB;
14'd14259:data <=32'h001BFFBC;14'd14260:data <=32'h000FFFAF;14'd14261:data <=32'hFFFEFFA4;
14'd14262:data <=32'hFFEAFF9F;14'd14263:data <=32'hFFD3FFA0;14'd14264:data <=32'hFFBEFFA8;
14'd14265:data <=32'hFFACFFB5;14'd14266:data <=32'hFF9FFFC6;14'd14267:data <=32'hFF96FFD8;
14'd14268:data <=32'hFF92FFEB;14'd14269:data <=32'hFF91FFFD;14'd14270:data <=32'hFF93000E;
14'd14271:data <=32'hFF98001F;14'd14272:data <=32'hFF93001C;14'd14273:data <=32'hFF920032;
14'd14274:data <=32'hFF940040;14'd14275:data <=32'hFF950028;14'd14276:data <=32'hFFAF0023;
14'd14277:data <=32'hFFB3002C;14'd14278:data <=32'hFFB80035;14'd14279:data <=32'hFFBD003D;
14'd14280:data <=32'hFFC40047;14'd14281:data <=32'hFFCB0051;14'd14282:data <=32'hFFD5005B;
14'd14283:data <=32'hFFE40064;14'd14284:data <=32'hFFF6006A;14'd14285:data <=32'h000B006B;
14'd14286:data <=32'h00200066;14'd14287:data <=32'h0032005B;14'd14288:data <=32'h0040004C;
14'd14289:data <=32'h004A003A;14'd14290:data <=32'h004D0027;14'd14291:data <=32'h004D0016;
14'd14292:data <=32'h00480007;14'd14293:data <=32'h0041FFFA;14'd14294:data <=32'h0038FFF0;
14'd14295:data <=32'h002DFFE9;14'd14296:data <=32'h0020FFE5;14'd14297:data <=32'h0014FFE5;
14'd14298:data <=32'h0008FFE8;14'd14299:data <=32'hFFFFFFF0;14'd14300:data <=32'hFFFAFFFA;
14'd14301:data <=32'hFFF90005;14'd14302:data <=32'hFFFD000F;14'd14303:data <=32'h00040016;
14'd14304:data <=32'h000E0019;14'd14305:data <=32'h00170019;14'd14306:data <=32'h001F0014;
14'd14307:data <=32'h0025000E;14'd14308:data <=32'h00270008;14'd14309:data <=32'h00270002;
14'd14310:data <=32'h0027FFFD;14'd14311:data <=32'h0026FFF9;14'd14312:data <=32'h0025FFF6;
14'd14313:data <=32'h0024FFF4;14'd14314:data <=32'h0023FFF1;14'd14315:data <=32'h0023FFEE;
14'd14316:data <=32'h0023FFEB;14'd14317:data <=32'h0022FFE8;14'd14318:data <=32'h0021FFE6;
14'd14319:data <=32'h0020FFE3;14'd14320:data <=32'h0021FFDF;14'd14321:data <=32'h0021FFDB;
14'd14322:data <=32'h001FFFD5;14'd14323:data <=32'h001DFFCE;14'd14324:data <=32'h0018FFC6;
14'd14325:data <=32'h0010FFBF;14'd14326:data <=32'h0006FFBA;14'd14327:data <=32'hFFFAFFB9;
14'd14328:data <=32'hFFEFFFBB;14'd14329:data <=32'hFFE5FFC0;14'd14330:data <=32'hFFDEFFC6;
14'd14331:data <=32'hFFDAFFCC;14'd14332:data <=32'hFFD8FFD1;14'd14333:data <=32'hFFD7FFD4;
14'd14334:data <=32'hFFD4FFD6;14'd14335:data <=32'hFFD0FFD6;14'd14336:data <=32'hFF99FFBD;
14'd14337:data <=32'hFF87FFCF;14'd14338:data <=32'hFF84FFE3;14'd14339:data <=32'hFFBFFFD8;
14'd14340:data <=32'hFFCBFFCB;14'd14341:data <=32'hFFBFFFCE;14'd14342:data <=32'hFFB2FFD3;
14'd14343:data <=32'hFFA5FFDE;14'd14344:data <=32'hFF99FFEC;14'd14345:data <=32'hFF90FFFF;
14'd14346:data <=32'hFF8C0015;14'd14347:data <=32'hFF8E002E;14'd14348:data <=32'hFF980046;
14'd14349:data <=32'hFFA9005B;14'd14350:data <=32'hFFBF006B;14'd14351:data <=32'hFFD80073;
14'd14352:data <=32'hFFF10073;14'd14353:data <=32'h0008006E;14'd14354:data <=32'h001C0064;
14'd14355:data <=32'h002B0056;14'd14356:data <=32'h00360047;14'd14357:data <=32'h003D0037;
14'd14358:data <=32'h00400026;14'd14359:data <=32'h003F0016;14'd14360:data <=32'h003A0007;
14'd14361:data <=32'h0032FFFA;14'd14362:data <=32'h0027FFF2;14'd14363:data <=32'h001AFFED;
14'd14364:data <=32'h000EFFED;14'd14365:data <=32'h0004FFF1;14'd14366:data <=32'hFFFCFFF8;
14'd14367:data <=32'hFFF80000;14'd14368:data <=32'hFFF80008;14'd14369:data <=32'hFFF9000E;
14'd14370:data <=32'hFFFC0013;14'd14371:data <=32'hFFFE0017;14'd14372:data <=32'h0000001A;
14'd14373:data <=32'h0003001E;14'd14374:data <=32'h00080023;14'd14375:data <=32'h000D0027;
14'd14376:data <=32'h0015002A;14'd14377:data <=32'h001F002B;14'd14378:data <=32'h002A002B;
14'd14379:data <=32'h00350026;14'd14380:data <=32'h003F001D;14'd14381:data <=32'h00470013;
14'd14382:data <=32'h004D0007;14'd14383:data <=32'h0050FFF9;14'd14384:data <=32'h004FFFEC;
14'd14385:data <=32'h004DFFDF;14'd14386:data <=32'h0048FFD2;14'd14387:data <=32'h0040FFC6;
14'd14388:data <=32'h0035FFBB;14'd14389:data <=32'h0028FFB3;14'd14390:data <=32'h0018FFAF;
14'd14391:data <=32'h0008FFAF;14'd14392:data <=32'hFFF9FFB4;14'd14393:data <=32'hFFEDFFBE;
14'd14394:data <=32'hFFE6FFCA;14'd14395:data <=32'hFFE5FFD5;14'd14396:data <=32'hFFE8FFDF;
14'd14397:data <=32'hFFEEFFE4;14'd14398:data <=32'hFFF5FFE5;14'd14399:data <=32'hFFFAFFE2;
14'd14400:data <=32'hFFF4FFAA;14'd14401:data <=32'hFFE3FFA5;14'd14402:data <=32'hFFD3FFAF;
14'd14403:data <=32'hFFE6FFDA;14'd14404:data <=32'hFFF8FFC7;14'd14405:data <=32'hFFF0FFC1;
14'd14406:data <=32'hFFE5FFBD;14'd14407:data <=32'hFFD9FFBC;14'd14408:data <=32'hFFCAFFBD;
14'd14409:data <=32'hFFBBFFC4;14'd14410:data <=32'hFFACFFCF;14'd14411:data <=32'hFFA1FFDF;
14'd14412:data <=32'hFF9BFFF3;14'd14413:data <=32'hFF9B0007;14'd14414:data <=32'hFFA0001A;
14'd14415:data <=32'hFFAA002A;14'd14416:data <=32'hFFB70035;14'd14417:data <=32'hFFC4003D;
14'd14418:data <=32'hFFD10041;14'd14419:data <=32'hFFDD0042;14'd14420:data <=32'hFFE80043;
14'd14421:data <=32'hFFF20042;14'd14422:data <=32'hFFFC0040;14'd14423:data <=32'h0005003B;
14'd14424:data <=32'h000E0036;14'd14425:data <=32'h0013002E;14'd14426:data <=32'h00170026;
14'd14427:data <=32'h0019001E;14'd14428:data <=32'h00180017;14'd14429:data <=32'h00160012;
14'd14430:data <=32'h0014000D;14'd14431:data <=32'h00120009;14'd14432:data <=32'h000F0005;
14'd14433:data <=32'h000C0002;14'd14434:data <=32'h0007FFFF;14'd14435:data <=32'h0001FFFC;
14'd14436:data <=32'hFFF9FFFD;14'd14437:data <=32'hFFF00000;14'd14438:data <=32'hFFE80008;
14'd14439:data <=32'hFFE30013;14'd14440:data <=32'hFFE10021;14'd14441:data <=32'hFFE5002F;
14'd14442:data <=32'hFFEE003C;14'd14443:data <=32'hFFFC0046;14'd14444:data <=32'h000C004C;
14'd14445:data <=32'h001D004E;14'd14446:data <=32'h002F004B;14'd14447:data <=32'h003F0043;
14'd14448:data <=32'h004D0039;14'd14449:data <=32'h0059002A;14'd14450:data <=32'h0062001A;
14'd14451:data <=32'h00670007;14'd14452:data <=32'h0067FFF3;14'd14453:data <=32'h0062FFDF;
14'd14454:data <=32'h0058FFCE;14'd14455:data <=32'h004AFFC0;14'd14456:data <=32'h0039FFB8;
14'd14457:data <=32'h0029FFB6;14'd14458:data <=32'h001AFFB8;14'd14459:data <=32'h000FFFBE;
14'd14460:data <=32'h0009FFC5;14'd14461:data <=32'h0006FFCB;14'd14462:data <=32'h0005FFCE;
14'd14463:data <=32'h0006FFCF;14'd14464:data <=32'h000FFFDE;14'd14465:data <=32'h0012FFD6;
14'd14466:data <=32'h000AFFCD;14'd14467:data <=32'hFFEFFFBE;14'd14468:data <=32'hFFFDFFB1;
14'd14469:data <=32'hFFF3FFB2;14'd14470:data <=32'hFFE9FFB4;14'd14471:data <=32'hFFE0FFB9;
14'd14472:data <=32'hFFD6FFBD;14'd14473:data <=32'hFFCDFFC4;14'd14474:data <=32'hFFC5FFCD;
14'd14475:data <=32'hFFBEFFD9;14'd14476:data <=32'hFFBBFFE5;14'd14477:data <=32'hFFBDFFF3;
14'd14478:data <=32'hFFC1FFFE;14'd14479:data <=32'hFFC90006;14'd14480:data <=32'hFFD1000A;
14'd14481:data <=32'hFFD8000A;14'd14482:data <=32'hFFDD0008;14'd14483:data <=32'hFFDF0006;
14'd14484:data <=32'hFFDD0005;14'd14485:data <=32'hFFDB0006;14'd14486:data <=32'hFFD90008;
14'd14487:data <=32'hFFD8000D;14'd14488:data <=32'hFFD80012;14'd14489:data <=32'hFFDA0017;
14'd14490:data <=32'hFFDD001C;14'd14491:data <=32'hFFE10020;14'd14492:data <=32'hFFE50024;
14'd14493:data <=32'hFFEB0027;14'd14494:data <=32'hFFF10029;14'd14495:data <=32'hFFF90029;
14'd14496:data <=32'h00010027;14'd14497:data <=32'h00090022;14'd14498:data <=32'h000E001A;
14'd14499:data <=32'h000F0010;14'd14500:data <=32'h000D0007;14'd14501:data <=32'h0007FFFE;
14'd14502:data <=32'hFFFCFFFA;14'd14503:data <=32'hFFF1FFFA;14'd14504:data <=32'hFFE7FFFF;
14'd14505:data <=32'hFFDF0008;14'd14506:data <=32'hFFDA0013;14'd14507:data <=32'hFFDA0020;
14'd14508:data <=32'hFFDD002C;14'd14509:data <=32'hFFE40036;14'd14510:data <=32'hFFED003F;
14'd14511:data <=32'hFFF70046;14'd14512:data <=32'h0003004A;14'd14513:data <=32'h0010004D;
14'd14514:data <=32'h001D004D;14'd14515:data <=32'h002C0049;14'd14516:data <=32'h00380043;
14'd14517:data <=32'h00440039;14'd14518:data <=32'h004C002D;14'd14519:data <=32'h00520021;
14'd14520:data <=32'h00540015;14'd14521:data <=32'h0054000B;14'd14522:data <=32'h00530002;
14'd14523:data <=32'h0053FFFA;14'd14524:data <=32'h0054FFF2;14'd14525:data <=32'h0055FFE8;
14'd14526:data <=32'h0055FFDD;14'd14527:data <=32'h0054FFD0;14'd14528:data <=32'h000CFFDF;
14'd14529:data <=32'h0011FFE2;14'd14530:data <=32'h001BFFDE;14'd14531:data <=32'h0041FFAF;
14'd14532:data <=32'h0047FF95;14'd14533:data <=32'h0031FF8C;14'd14534:data <=32'h001AFF88;
14'd14535:data <=32'h0003FF89;14'd14536:data <=32'hFFEEFF8E;14'd14537:data <=32'hFFDAFF98;
14'd14538:data <=32'hFFCAFFA5;14'd14539:data <=32'hFFBDFFB7;14'd14540:data <=32'hFFB5FFCB;
14'd14541:data <=32'hFFB4FFDF;14'd14542:data <=32'hFFB9FFF2;14'd14543:data <=32'hFFC30001;
14'd14544:data <=32'hFFD1000A;14'd14545:data <=32'hFFDF000D;14'd14546:data <=32'hFFEA000B;
14'd14547:data <=32'hFFF30005;14'd14548:data <=32'hFFF7FFFD;14'd14549:data <=32'hFFF7FFF7;
14'd14550:data <=32'hFFF4FFF1;14'd14551:data <=32'hFFEFFFEE;14'd14552:data <=32'hFFEBFFED;
14'd14553:data <=32'hFFE6FFED;14'd14554:data <=32'hFFE1FFEF;14'd14555:data <=32'hFFDCFFF2;
14'd14556:data <=32'hFFD8FFF6;14'd14557:data <=32'hFFD5FFFD;14'd14558:data <=32'hFFD40004;
14'd14559:data <=32'hFFD5000B;14'd14560:data <=32'hFFD90012;14'd14561:data <=32'hFFDF0016;
14'd14562:data <=32'hFFE60019;14'd14563:data <=32'hFFEC0018;14'd14564:data <=32'hFFF00016;
14'd14565:data <=32'hFFF30011;14'd14566:data <=32'hFFF2000E;14'd14567:data <=32'hFFF0000B;
14'd14568:data <=32'hFFED000C;14'd14569:data <=32'hFFEA000D;14'd14570:data <=32'hFFE80011;
14'd14571:data <=32'hFFE80014;14'd14572:data <=32'hFFE90017;14'd14573:data <=32'hFFEB001A;
14'd14574:data <=32'hFFEC001B;14'd14575:data <=32'hFFED001C;14'd14576:data <=32'hFFEC001E;
14'd14577:data <=32'hFFEB0021;14'd14578:data <=32'hFFEB0025;14'd14579:data <=32'hFFEB002B;
14'd14580:data <=32'hFFEE0031;14'd14581:data <=32'hFFF10037;14'd14582:data <=32'hFFF7003D;
14'd14583:data <=32'hFFFD0043;14'd14584:data <=32'h00050049;14'd14585:data <=32'h000E004E;
14'd14586:data <=32'h001A0054;14'd14587:data <=32'h00290057;14'd14588:data <=32'h003B0058;
14'd14589:data <=32'h004F0053;14'd14590:data <=32'h00640048;14'd14591:data <=32'h00770036;
14'd14592:data <=32'h0039FFFA;14'd14593:data <=32'h003EFFF8;14'd14594:data <=32'h0045FFFD;
14'd14595:data <=32'h0077000F;14'd14596:data <=32'h008DFFE8;14'd14597:data <=32'h0084FFCE;
14'd14598:data <=32'h0075FFB8;14'd14599:data <=32'h0062FFA6;14'd14600:data <=32'h004EFF98;
14'd14601:data <=32'h0036FF90;14'd14602:data <=32'h001EFF8D;14'd14603:data <=32'h0006FF90;
14'd14604:data <=32'hFFF1FF99;14'd14605:data <=32'hFFE0FFA7;14'd14606:data <=32'hFFD5FFB7;
14'd14607:data <=32'hFFD0FFC8;14'd14608:data <=32'hFFD1FFD8;14'd14609:data <=32'hFFD5FFE4;
14'd14610:data <=32'hFFDBFFEB;14'd14611:data <=32'hFFE1FFF0;14'd14612:data <=32'hFFE6FFF2;
14'd14613:data <=32'hFFE8FFF3;14'd14614:data <=32'hFFEAFFF4;14'd14615:data <=32'hFFEBFFF5;
14'd14616:data <=32'hFFEEFFF6;14'd14617:data <=32'hFFF0FFF7;14'd14618:data <=32'hFFF3FFF6;
14'd14619:data <=32'hFFF4FFF5;14'd14620:data <=32'hFFF5FFF2;14'd14621:data <=32'hFFF4FFF0;
14'd14622:data <=32'hFFF2FFEE;14'd14623:data <=32'hFFF0FFED;14'd14624:data <=32'hFFEDFFED;
14'd14625:data <=32'hFFEBFFED;14'd14626:data <=32'hFFE9FFED;14'd14627:data <=32'hFFE7FFED;
14'd14628:data <=32'hFFE3FFED;14'd14629:data <=32'hFFDFFFED;14'd14630:data <=32'hFFDAFFEF;
14'd14631:data <=32'hFFD3FFF3;14'd14632:data <=32'hFFCEFFFA;14'd14633:data <=32'hFFCB0003;
14'd14634:data <=32'hFFCB000D;14'd14635:data <=32'hFFCF0016;14'd14636:data <=32'hFFD6001D;
14'd14637:data <=32'hFFDF0022;14'd14638:data <=32'hFFE70022;14'd14639:data <=32'hFFEE0020;
14'd14640:data <=32'hFFF2001C;14'd14641:data <=32'hFFF40016;14'd14642:data <=32'hFFF30012;
14'd14643:data <=32'hFFEF0010;14'd14644:data <=32'hFFEA000E;14'd14645:data <=32'hFFE50010;
14'd14646:data <=32'hFFDF0014;14'd14647:data <=32'hFFDA001A;14'd14648:data <=32'hFFD50023;
14'd14649:data <=32'hFFD3002F;14'd14650:data <=32'hFFD4003E;14'd14651:data <=32'hFFDA004E;
14'd14652:data <=32'hFFE6005D;14'd14653:data <=32'hFFF7006B;14'd14654:data <=32'h000E0073;
14'd14655:data <=32'h00280075;14'd14656:data <=32'h001F0050;14'd14657:data <=32'h00330054;
14'd14658:data <=32'h003D0054;14'd14659:data <=32'h00360056;14'd14660:data <=32'h005A003D;
14'd14661:data <=32'h0061002E;14'd14662:data <=32'h0064001D;14'd14663:data <=32'h0065000E;
14'd14664:data <=32'h0063FFFF;14'd14665:data <=32'h0060FFF0;14'd14666:data <=32'h0059FFE2;
14'd14667:data <=32'h0051FFD6;14'd14668:data <=32'h0046FFCE;14'd14669:data <=32'h003BFFC8;
14'd14670:data <=32'h0030FFC5;14'd14671:data <=32'h0028FFC4;14'd14672:data <=32'h0020FFC4;
14'd14673:data <=32'h001AFFC3;14'd14674:data <=32'h0014FFC2;14'd14675:data <=32'h000CFFBF;
14'd14676:data <=32'h0003FFBE;14'd14677:data <=32'hFFF8FFC0;14'd14678:data <=32'hFFEDFFC4;
14'd14679:data <=32'hFFE4FFCB;14'd14680:data <=32'hFFDCFFD6;14'd14681:data <=32'hFFDAFFE2;
14'd14682:data <=32'hFFDAFFED;14'd14683:data <=32'hFFDFFFF7;14'd14684:data <=32'hFFE6FFFE;
14'd14685:data <=32'hFFED0002;14'd14686:data <=32'hFFF50004;14'd14687:data <=32'hFFFD0003;
14'd14688:data <=32'h00040000;14'd14689:data <=32'h0009FFFB;14'd14690:data <=32'h000DFFF4;
14'd14691:data <=32'h000FFFEC;14'd14692:data <=32'h000EFFE2;14'd14693:data <=32'h0009FFD8;
14'd14694:data <=32'h0000FFD0;14'd14695:data <=32'hFFF5FFCA;14'd14696:data <=32'hFFE8FFCA;
14'd14697:data <=32'hFFDBFFCD;14'd14698:data <=32'hFFCFFFD5;14'd14699:data <=32'hFFC7FFE0;
14'd14700:data <=32'hFFC4FFEC;14'd14701:data <=32'hFFC4FFF7;14'd14702:data <=32'hFFC70000;
14'd14703:data <=32'hFFCB0006;14'd14704:data <=32'hFFCF000A;14'd14705:data <=32'hFFD3000C;
14'd14706:data <=32'hFFD5000D;14'd14707:data <=32'hFFD6000E;14'd14708:data <=32'hFFD60010;
14'd14709:data <=32'hFFD60012;14'd14710:data <=32'hFFD50014;14'd14711:data <=32'hFFD40018;
14'd14712:data <=32'hFFD3001C;14'd14713:data <=32'hFFD10021;14'd14714:data <=32'hFFD00029;
14'd14715:data <=32'hFFD00033;14'd14716:data <=32'hFFD4003E;14'd14717:data <=32'hFFDB0049;
14'd14718:data <=32'hFFE70053;14'd14719:data <=32'hFFF6005A;14'd14720:data <=32'hFFC0004D;
14'd14721:data <=32'hFFCD0067;14'd14722:data <=32'hFFE20072;14'd14723:data <=32'h00060045;
14'd14724:data <=32'h00230034;14'd14725:data <=32'h0024002D;14'd14726:data <=32'h00230028;
14'd14727:data <=32'h00210026;14'd14728:data <=32'h00210025;14'd14729:data <=32'h00230026;
14'd14730:data <=32'h00270025;14'd14731:data <=32'h002B0024;14'd14732:data <=32'h00300022;
14'd14733:data <=32'h00350020;14'd14734:data <=32'h003B001C;14'd14735:data <=32'h00420017;
14'd14736:data <=32'h0049000F;14'd14737:data <=32'h004F0005;14'd14738:data <=32'h0054FFF6;
14'd14739:data <=32'h0054FFE6;14'd14740:data <=32'h004FFFD5;14'd14741:data <=32'h0044FFC5;
14'd14742:data <=32'h0035FFBA;14'd14743:data <=32'h0023FFB3;14'd14744:data <=32'h0010FFB3;
14'd14745:data <=32'hFFFFFFB8;14'd14746:data <=32'hFFF2FFC0;14'd14747:data <=32'hFFE8FFCC;
14'd14748:data <=32'hFFE3FFD8;14'd14749:data <=32'hFFE1FFE4;14'd14750:data <=32'hFFE2FFEF;
14'd14751:data <=32'hFFE7FFF9;14'd14752:data <=32'hFFEC0001;14'd14753:data <=32'hFFF50007;
14'd14754:data <=32'hFFFF000A;14'd14755:data <=32'h00090009;14'd14756:data <=32'h00130004;
14'd14757:data <=32'h001AFFFD;14'd14758:data <=32'h001EFFF2;14'd14759:data <=32'h001FFFE7;
14'd14760:data <=32'h001CFFDD;14'd14761:data <=32'h0015FFD4;14'd14762:data <=32'h000DFFCE;
14'd14763:data <=32'h0006FFCA;14'd14764:data <=32'hFFFEFFC9;14'd14765:data <=32'hFFF7FFC8;
14'd14766:data <=32'hFFF0FFC7;14'd14767:data <=32'hFFEAFFC6;14'd14768:data <=32'hFFE1FFC5;
14'd14769:data <=32'hFFD8FFC5;14'd14770:data <=32'hFFCDFFC7;14'd14771:data <=32'hFFC1FFCC;
14'd14772:data <=32'hFFB5FFD5;14'd14773:data <=32'hFFACFFE0;14'd14774:data <=32'hFFA5FFEE;
14'd14775:data <=32'hFFA1FFFC;14'd14776:data <=32'hFFA1000C;14'd14777:data <=32'hFFA2001B;
14'd14778:data <=32'hFFA6002A;14'd14779:data <=32'hFFAD0038;14'd14780:data <=32'hFFB70045;
14'd14781:data <=32'hFFC40051;14'd14782:data <=32'hFFD4005A;14'd14783:data <=32'hFFE7005E;
14'd14784:data <=32'hFFAE000B;14'd14785:data <=32'hFFA70023;14'd14786:data <=32'hFFAF003F;
14'd14787:data <=32'hFFFA0052;14'd14788:data <=32'h001B003D;14'd14789:data <=32'h001D002F;
14'd14790:data <=32'h001A0024;14'd14791:data <=32'h0014001D;14'd14792:data <=32'h000E001A;
14'd14793:data <=32'h0009001A;14'd14794:data <=32'h0005001C;14'd14795:data <=32'h00040021;
14'd14796:data <=32'h00040025;14'd14797:data <=32'h0006002B;14'd14798:data <=32'h000A0030;
14'd14799:data <=32'h00120036;14'd14800:data <=32'h001C0038;14'd14801:data <=32'h00290038;
14'd14802:data <=32'h00370033;14'd14803:data <=32'h00430029;14'd14804:data <=32'h004C001B;
14'd14805:data <=32'h004F000B;14'd14806:data <=32'h004EFFFB;14'd14807:data <=32'h0048FFEC;
14'd14808:data <=32'h003FFFE1;14'd14809:data <=32'h0034FFDA;14'd14810:data <=32'h0029FFD6;
14'd14811:data <=32'h001FFFD5;14'd14812:data <=32'h0017FFD5;14'd14813:data <=32'h000FFFD7;
14'd14814:data <=32'h0008FFDA;14'd14815:data <=32'h0002FFDE;14'd14816:data <=32'hFFFEFFE3;
14'd14817:data <=32'hFFFAFFE9;14'd14818:data <=32'hFFF8FFEF;14'd14819:data <=32'hFFFAFFF6;
14'd14820:data <=32'hFFFDFFFC;14'd14821:data <=32'h00010000;14'd14822:data <=32'h00070002;
14'd14823:data <=32'h000C0002;14'd14824:data <=32'h00110001;14'd14825:data <=32'h0016FFFF;
14'd14826:data <=32'h001BFFFD;14'd14827:data <=32'h001FFFF9;14'd14828:data <=32'h0025FFF5;
14'd14829:data <=32'h002BFFED;14'd14830:data <=32'h002FFFE3;14'd14831:data <=32'h0032FFD6;
14'd14832:data <=32'h0031FFC6;14'd14833:data <=32'h002AFFB6;14'd14834:data <=32'h001DFFA5;
14'd14835:data <=32'h000BFF99;14'd14836:data <=32'hFFF6FF92;14'd14837:data <=32'hFFDDFF91;
14'd14838:data <=32'hFFC6FF96;14'd14839:data <=32'hFFB0FFA0;14'd14840:data <=32'hFF9EFFAF;
14'd14841:data <=32'hFF8EFFC2;14'd14842:data <=32'hFF84FFD8;14'd14843:data <=32'hFF7EFFF1;
14'd14844:data <=32'hFF7D000A;14'd14845:data <=32'hFF830023;14'd14846:data <=32'hFF8F003A;
14'd14847:data <=32'hFFA1004D;14'd14848:data <=32'hFFBC0002;14'd14849:data <=32'hFFB3000F;
14'd14850:data <=32'hFFAB0022;14'd14851:data <=32'hFFB0004E;14'd14852:data <=32'hFFD90046;
14'd14853:data <=32'hFFE40042;14'd14854:data <=32'hFFEB003E;14'd14855:data <=32'hFFEF003A;
14'd14856:data <=32'hFFF30038;14'd14857:data <=32'hFFF70037;14'd14858:data <=32'hFFFA0036;
14'd14859:data <=32'hFFFF0035;14'd14860:data <=32'h00020034;14'd14861:data <=32'h00060032;
14'd14862:data <=32'h00090031;14'd14863:data <=32'h000D0031;14'd14864:data <=32'h00110031;
14'd14865:data <=32'h00160031;14'd14866:data <=32'h001D002E;14'd14867:data <=32'h00230029;
14'd14868:data <=32'h00280022;14'd14869:data <=32'h002B001A;14'd14870:data <=32'h002B0012;
14'd14871:data <=32'h0028000B;14'd14872:data <=32'h00240007;14'd14873:data <=32'h001F0005;
14'd14874:data <=32'h001C0005;14'd14875:data <=32'h001B0007;14'd14876:data <=32'h001C0007;
14'd14877:data <=32'h001E0007;14'd14878:data <=32'h00200005;14'd14879:data <=32'h00220001;
14'd14880:data <=32'h0022FFFC;14'd14881:data <=32'h0021FFF8;14'd14882:data <=32'h001EFFF4;
14'd14883:data <=32'h001AFFF2;14'd14884:data <=32'h0017FFF1;14'd14885:data <=32'h0013FFF0;
14'd14886:data <=32'h000FFFF1;14'd14887:data <=32'h000DFFF3;14'd14888:data <=32'h0009FFF5;
14'd14889:data <=32'h0008FFFA;14'd14890:data <=32'h0008FFFF;14'd14891:data <=32'h000A0005;
14'd14892:data <=32'h0010000B;14'd14893:data <=32'h0019000E;14'd14894:data <=32'h0025000F;
14'd14895:data <=32'h0032000A;14'd14896:data <=32'h003E0000;14'd14897:data <=32'h0047FFF0;
14'd14898:data <=32'h004BFFDE;14'd14899:data <=32'h0049FFCA;14'd14900:data <=32'h0040FFB7;
14'd14901:data <=32'h0033FFA6;14'd14902:data <=32'h0022FF9A;14'd14903:data <=32'h000FFF92;
14'd14904:data <=32'hFFFAFF8F;14'd14905:data <=32'hFFE6FF8F;14'd14906:data <=32'hFFD2FF94;
14'd14907:data <=32'hFFBFFF9D;14'd14908:data <=32'hFFAEFFAA;14'd14909:data <=32'hFFA0FFBB;
14'd14910:data <=32'hFF97FFCE;14'd14911:data <=32'hFF93FFE3;14'd14912:data <=32'hFF9DFFE4;
14'd14913:data <=32'hFF95FFF4;14'd14914:data <=32'hFF91FFFD;14'd14915:data <=32'hFF93FFE8;
14'd14916:data <=32'hFFABFFEB;14'd14917:data <=32'hFFA7FFF4;14'd14918:data <=32'hFFA3FFFE;
14'd14919:data <=32'hFFA0000A;14'd14920:data <=32'hFFA00019;14'd14921:data <=32'hFFA3002A;
14'd14922:data <=32'hFFAB003A;14'd14923:data <=32'hFFB70048;14'd14924:data <=32'hFFC50052;
14'd14925:data <=32'hFFD60059;14'd14926:data <=32'hFFE7005B;14'd14927:data <=32'hFFF7005A;
14'd14928:data <=32'h00060056;14'd14929:data <=32'h00140050;14'd14930:data <=32'h00200047;
14'd14931:data <=32'h002A003A;14'd14932:data <=32'h0031002C;14'd14933:data <=32'h0032001D;
14'd14934:data <=32'h002F000E;14'd14935:data <=32'h00280002;14'd14936:data <=32'h001DFFFB;
14'd14937:data <=32'h0011FFF8;14'd14938:data <=32'h0006FFFA;14'd14939:data <=32'hFFFE0000;
14'd14940:data <=32'hFFFA0009;14'd14941:data <=32'hFFFA0011;14'd14942:data <=32'hFFFD0018;
14'd14943:data <=32'h0002001C;14'd14944:data <=32'h0008001E;14'd14945:data <=32'h000E001F;
14'd14946:data <=32'h0013001E;14'd14947:data <=32'h0018001C;14'd14948:data <=32'h001C0019;
14'd14949:data <=32'h001F0015;14'd14950:data <=32'h00210011;14'd14951:data <=32'h0023000D;
14'd14952:data <=32'h00220008;14'd14953:data <=32'h00210005;14'd14954:data <=32'h001E0003;
14'd14955:data <=32'h001B0003;14'd14956:data <=32'h001B0005;14'd14957:data <=32'h001C0008;
14'd14958:data <=32'h0020000B;14'd14959:data <=32'h0027000B;14'd14960:data <=32'h002E0008;
14'd14961:data <=32'h00360002;14'd14962:data <=32'h003BFFF9;14'd14963:data <=32'h003DFFEE;
14'd14964:data <=32'h003CFFE3;14'd14965:data <=32'h0038FFD9;14'd14966:data <=32'h0032FFD1;
14'd14967:data <=32'h002CFFCB;14'd14968:data <=32'h0025FFC6;14'd14969:data <=32'h001FFFC2;
14'd14970:data <=32'h0018FFBE;14'd14971:data <=32'h0012FFBA;14'd14972:data <=32'h000AFFB7;
14'd14973:data <=32'h0001FFB5;14'd14974:data <=32'hFFF9FFB4;14'd14975:data <=32'hFFF0FFB5;
14'd14976:data <=32'hFFC6FF98;14'd14977:data <=32'hFFB2FFA1;14'd14978:data <=32'hFFADFFAE;
14'd14979:data <=32'hFFE6FFB0;14'd14980:data <=32'hFFF4FFA4;14'd14981:data <=32'hFFE3FF9E;
14'd14982:data <=32'hFFCFFF9E;14'd14983:data <=32'hFFB9FFA2;14'd14984:data <=32'hFFA3FFAE;
14'd14985:data <=32'hFF91FFC1;14'd14986:data <=32'hFF85FFD8;14'd14987:data <=32'hFF80FFF2;
14'd14988:data <=32'hFF81000C;14'd14989:data <=32'hFF890024;14'd14990:data <=32'hFF950038;
14'd14991:data <=32'hFFA50049;14'd14992:data <=32'hFFB80056;14'd14993:data <=32'hFFCC005E;
14'd14994:data <=32'hFFE20061;14'd14995:data <=32'hFFF7005F;14'd14996:data <=32'h000B0056;
14'd14997:data <=32'h001B004A;14'd14998:data <=32'h00250039;14'd14999:data <=32'h002A0027;
14'd15000:data <=32'h00290017;14'd15001:data <=32'h0022000A;14'd15002:data <=32'h00190001;
14'd15003:data <=32'h000FFFFC;14'd15004:data <=32'h0006FFFC;14'd15005:data <=32'hFFFFFFFD;
14'd15006:data <=32'hFFFA0000;14'd15007:data <=32'hFFF60004;14'd15008:data <=32'hFFF30008;
14'd15009:data <=32'hFFF1000C;14'd15010:data <=32'hFFEF0011;14'd15011:data <=32'hFFEE0016;
14'd15012:data <=32'hFFEF001C;14'd15013:data <=32'hFFF10023;14'd15014:data <=32'hFFF50029;
14'd15015:data <=32'hFFFB002E;14'd15016:data <=32'h00020032;14'd15017:data <=32'h000A0034;
14'd15018:data <=32'h00120034;14'd15019:data <=32'h001A0034;14'd15020:data <=32'h00220032;
14'd15021:data <=32'h002A0030;14'd15022:data <=32'h0033002D;14'd15023:data <=32'h003C0026;
14'd15024:data <=32'h0045001D;14'd15025:data <=32'h004B0012;14'd15026:data <=32'h004E0003;
14'd15027:data <=32'h004DFFF5;14'd15028:data <=32'h0047FFE7;14'd15029:data <=32'h003EFFDD;
14'd15030:data <=32'h0033FFD6;14'd15031:data <=32'h0028FFD4;14'd15032:data <=32'h001FFFD6;
14'd15033:data <=32'h0018FFD9;14'd15034:data <=32'h0014FFDE;14'd15035:data <=32'h0014FFE2;
14'd15036:data <=32'h0015FFE4;14'd15037:data <=32'h0018FFE5;14'd15038:data <=32'h001BFFE5;
14'd15039:data <=32'h001FFFE2;14'd15040:data <=32'h0025FFAD;14'd15041:data <=32'h001AFFA3;
14'd15042:data <=32'h000CFFA6;14'd15043:data <=32'h0017FFD4;14'd15044:data <=32'h0031FFC3;
14'd15045:data <=32'h002AFFB3;14'd15046:data <=32'h001DFFA5;14'd15047:data <=32'h000CFF9A;
14'd15048:data <=32'hFFF7FF95;14'd15049:data <=32'hFFE0FF96;14'd15050:data <=32'hFFCBFF9E;
14'd15051:data <=32'hFFBAFFAB;14'd15052:data <=32'hFFADFFBA;14'd15053:data <=32'hFFA4FFCC;
14'd15054:data <=32'hFFA0FFDD;14'd15055:data <=32'hFF9EFFEE;14'd15056:data <=32'hFFA0FFFF;
14'd15057:data <=32'hFFA5000F;14'd15058:data <=32'hFFAD001E;14'd15059:data <=32'hFFB80029;
14'd15060:data <=32'hFFC50032;14'd15061:data <=32'hFFD30036;14'd15062:data <=32'hFFE00037;
14'd15063:data <=32'hFFEC0034;14'd15064:data <=32'hFFF5002F;14'd15065:data <=32'hFFFB0029;
14'd15066:data <=32'hFFFF0024;14'd15067:data <=32'h00010020;14'd15068:data <=32'h0004001C;
14'd15069:data <=32'h00060018;14'd15070:data <=32'h00090014;14'd15071:data <=32'h000A000E;
14'd15072:data <=32'h000A0007;14'd15073:data <=32'h00070000;14'd15074:data <=32'h0001FFFA;
14'd15075:data <=32'hFFF8FFF6;14'd15076:data <=32'hFFEEFFF6;14'd15077:data <=32'hFFE4FFF9;
14'd15078:data <=32'hFFDB0000;14'd15079:data <=32'hFFD5000A;14'd15080:data <=32'hFFD20015;
14'd15081:data <=32'hFFD10022;14'd15082:data <=32'hFFD4002E;14'd15083:data <=32'hFFDA003B;
14'd15084:data <=32'hFFE20047;14'd15085:data <=32'hFFEF0051;14'd15086:data <=32'hFFFE0058;
14'd15087:data <=32'h0011005C;14'd15088:data <=32'h0024005A;14'd15089:data <=32'h00370053;
14'd15090:data <=32'h00470046;14'd15091:data <=32'h00530035;14'd15092:data <=32'h00590022;
14'd15093:data <=32'h00590010;14'd15094:data <=32'h0055FFFF;14'd15095:data <=32'h004CFFF3;
14'd15096:data <=32'h0043FFEB;14'd15097:data <=32'h0039FFE7;14'd15098:data <=32'h0031FFE5;
14'd15099:data <=32'h002BFFE6;14'd15100:data <=32'h0027FFE7;14'd15101:data <=32'h0025FFE8;
14'd15102:data <=32'h0024FFE9;14'd15103:data <=32'h0025FFEA;14'd15104:data <=32'h0028FFF6;
14'd15105:data <=32'h0030FFF2;14'd15106:data <=32'h0030FFE9;14'd15107:data <=32'h001EFFD7;
14'd15108:data <=32'h0036FFCD;14'd15109:data <=32'h0031FFC4;14'd15110:data <=32'h0029FFBA;
14'd15111:data <=32'h001EFFB3;14'd15112:data <=32'h0010FFAE;14'd15113:data <=32'h0001FFAE;
14'd15114:data <=32'hFFF4FFB3;14'd15115:data <=32'hFFE9FFBA;14'd15116:data <=32'hFFE2FFC3;
14'd15117:data <=32'hFFDEFFCB;14'd15118:data <=32'hFFDDFFD2;14'd15119:data <=32'hFFDCFFD8;
14'd15120:data <=32'hFFDBFFDC;14'd15121:data <=32'hFFDAFFDF;14'd15122:data <=32'hFFD8FFE3;
14'd15123:data <=32'hFFD6FFE7;14'd15124:data <=32'hFFD5FFEB;14'd15125:data <=32'hFFD5FFEF;
14'd15126:data <=32'hFFD5FFF2;14'd15127:data <=32'hFFD3FFF5;14'd15128:data <=32'hFFD2FFF8;
14'd15129:data <=32'hFFD0FFFD;14'd15130:data <=32'hFFCF0003;14'd15131:data <=32'hFFCF000B;
14'd15132:data <=32'hFFD10014;14'd15133:data <=32'hFFD8001C;14'd15134:data <=32'hFFE10022;
14'd15135:data <=32'hFFEC0024;14'd15136:data <=32'hFFF70022;14'd15137:data <=32'h0001001C;
14'd15138:data <=32'h00060013;14'd15139:data <=32'h00080008;14'd15140:data <=32'h0006FFFF;
14'd15141:data <=32'h0000FFF6;14'd15142:data <=32'hFFF8FFF1;14'd15143:data <=32'hFFEEFFEF;
14'd15144:data <=32'hFFE4FFEF;14'd15145:data <=32'hFFDAFFF3;14'd15146:data <=32'hFFD1FFFA;
14'd15147:data <=32'hFFC90003;14'd15148:data <=32'hFFC4000F;14'd15149:data <=32'hFFC2001D;
14'd15150:data <=32'hFFC3002C;14'd15151:data <=32'hFFCA003B;14'd15152:data <=32'hFFD40048;
14'd15153:data <=32'hFFE10052;14'd15154:data <=32'hFFF10058;14'd15155:data <=32'h00020058;
14'd15156:data <=32'h00100055;14'd15157:data <=32'h001C0050;14'd15158:data <=32'h00250049;
14'd15159:data <=32'h002C0043;14'd15160:data <=32'h0032003D;14'd15161:data <=32'h00370039;
14'd15162:data <=32'h003E0034;14'd15163:data <=32'h0045002E;14'd15164:data <=32'h004C0027;
14'd15165:data <=32'h0053001D;14'd15166:data <=32'h00570011;14'd15167:data <=32'h005A0005;
14'd15168:data <=32'h000FFFFC;14'd15169:data <=32'h00140006;14'd15170:data <=32'h0023000A;
14'd15171:data <=32'h0059FFEA;14'd15172:data <=32'h006EFFD6;14'd15173:data <=32'h0064FFC4;
14'd15174:data <=32'h0055FFB3;14'd15175:data <=32'h0042FFA6;14'd15176:data <=32'h002DFF9F;
14'd15177:data <=32'h0016FF9F;14'd15178:data <=32'h0001FFA5;14'd15179:data <=32'hFFF1FFB1;
14'd15180:data <=32'hFFE6FFBF;14'd15181:data <=32'hFFE2FFCE;14'd15182:data <=32'hFFE2FFDB;
14'd15183:data <=32'hFFE6FFE6;14'd15184:data <=32'hFFECFFEC;14'd15185:data <=32'hFFF2FFEF;
14'd15186:data <=32'hFFF8FFF0;14'd15187:data <=32'hFFFCFFEF;14'd15188:data <=32'hFFFFFFEB;
14'd15189:data <=32'h0001FFE7;14'd15190:data <=32'h0001FFE3;14'd15191:data <=32'hFFFFFFDD;
14'd15192:data <=32'hFFFAFFD8;14'd15193:data <=32'hFFF2FFD4;14'd15194:data <=32'hFFE8FFD4;
14'd15195:data <=32'hFFDFFFD8;14'd15196:data <=32'hFFD6FFDE;14'd15197:data <=32'hFFD1FFE8;
14'd15198:data <=32'hFFCFFFF3;14'd15199:data <=32'hFFD2FFFD;14'd15200:data <=32'hFFD80005;
14'd15201:data <=32'hFFDF0009;14'd15202:data <=32'hFFE6000A;14'd15203:data <=32'hFFEB0009;
14'd15204:data <=32'hFFEF0006;14'd15205:data <=32'hFFF00003;14'd15206:data <=32'hFFF10000;
14'd15207:data <=32'hFFF0FFFE;14'd15208:data <=32'hFFEFFFFC;14'd15209:data <=32'hFFEDFFFB;
14'd15210:data <=32'hFFEAFFF9;14'd15211:data <=32'hFFE7FFF8;14'd15212:data <=32'hFFE3FFF8;
14'd15213:data <=32'hFFDEFFF9;14'd15214:data <=32'hFFD8FFFC;14'd15215:data <=32'hFFD40001;
14'd15216:data <=32'hFFD00007;14'd15217:data <=32'hFFCE000D;14'd15218:data <=32'hFFCE0014;
14'd15219:data <=32'hFFCE001A;14'd15220:data <=32'hFFCE0020;14'd15221:data <=32'hFFCD0026;
14'd15222:data <=32'hFFCD002F;14'd15223:data <=32'hFFCD0039;14'd15224:data <=32'hFFCF0046;
14'd15225:data <=32'hFFD60054;14'd15226:data <=32'hFFE20063;14'd15227:data <=32'hFFF3006F;
14'd15228:data <=32'h00080076;14'd15229:data <=32'h001F0078;14'd15230:data <=32'h00370074;
14'd15231:data <=32'h004E006A;14'd15232:data <=32'h00220014;14'd15233:data <=32'h0024001B;
14'd15234:data <=32'h0029002A;14'd15235:data <=32'h005B0050;14'd15236:data <=32'h00830038;
14'd15237:data <=32'h008A001D;14'd15238:data <=32'h00890000;14'd15239:data <=32'h0082FFE5;
14'd15240:data <=32'h0074FFCD;14'd15241:data <=32'h0060FFBB;14'd15242:data <=32'h0049FFB0;
14'd15243:data <=32'h0033FFAD;14'd15244:data <=32'h001FFFB0;14'd15245:data <=32'h000FFFB7;
14'd15246:data <=32'h0004FFC1;14'd15247:data <=32'hFFFEFFCB;14'd15248:data <=32'hFFFBFFD3;
14'd15249:data <=32'hFFF9FFDA;14'd15250:data <=32'hFFF8FFE0;14'd15251:data <=32'hFFF9FFE5;
14'd15252:data <=32'hFFFBFFE9;14'd15253:data <=32'hFFFDFFEC;14'd15254:data <=32'h0000FFEE;
14'd15255:data <=32'h0004FFED;14'd15256:data <=32'h0006FFEB;14'd15257:data <=32'h0006FFE7;
14'd15258:data <=32'h0004FFE3;14'd15259:data <=32'h0001FFE1;14'd15260:data <=32'hFFFDFFE0;
14'd15261:data <=32'hFFF9FFE1;14'd15262:data <=32'hFFF7FFE4;14'd15263:data <=32'hFFF6FFE6;
14'd15264:data <=32'hFFF6FFE7;14'd15265:data <=32'hFFF7FFE6;14'd15266:data <=32'hFFF7FFE4;
14'd15267:data <=32'hFFF5FFE2;14'd15268:data <=32'hFFF1FFDF;14'd15269:data <=32'hFFEBFFDF;
14'd15270:data <=32'hFFE5FFE0;14'd15271:data <=32'hFFDFFFE4;14'd15272:data <=32'hFFDBFFEA;
14'd15273:data <=32'hFFD9FFF0;14'd15274:data <=32'hFFDAFFF6;14'd15275:data <=32'hFFDCFFFB;
14'd15276:data <=32'hFFDFFFFF;14'd15277:data <=32'hFFE20001;14'd15278:data <=32'hFFE50001;
14'd15279:data <=32'hFFE70000;14'd15280:data <=32'hFFE9FFFF;14'd15281:data <=32'hFFEAFFFC;
14'd15282:data <=32'hFFE9FFF9;14'd15283:data <=32'hFFE7FFF5;14'd15284:data <=32'hFFE1FFF0;
14'd15285:data <=32'hFFD9FFED;14'd15286:data <=32'hFFCDFFED;14'd15287:data <=32'hFFBFFFF2;
14'd15288:data <=32'hFFB2FFFD;14'd15289:data <=32'hFFA7000D;14'd15290:data <=32'hFFA20022;
14'd15291:data <=32'hFFA2003A;14'd15292:data <=32'hFFAB0051;14'd15293:data <=32'hFFB90066;
14'd15294:data <=32'hFFCE0076;14'd15295:data <=32'hFFE50081;14'd15296:data <=32'hFFF1004E;
14'd15297:data <=32'hFFFA005B;14'd15298:data <=32'hFFFD0065;14'd15299:data <=32'hFFF60074;
14'd15300:data <=32'h00260070;14'd15301:data <=32'h00390066;14'd15302:data <=32'h00480059;
14'd15303:data <=32'h00540048;14'd15304:data <=32'h005B0036;14'd15305:data <=32'h005D0024;
14'd15306:data <=32'h005A0014;14'd15307:data <=32'h00550007;14'd15308:data <=32'h0050FFFE;
14'd15309:data <=32'h004BFFF7;14'd15310:data <=32'h0047FFF1;14'd15311:data <=32'h0043FFEB;
14'd15312:data <=32'h0040FFE4;14'd15313:data <=32'h003BFFDC;14'd15314:data <=32'h0034FFD5;
14'd15315:data <=32'h002BFFCF;14'd15316:data <=32'h0021FFCC;14'd15317:data <=32'h0017FFCC;
14'd15318:data <=32'h000DFFCD;14'd15319:data <=32'h0005FFD1;14'd15320:data <=32'hFFFFFFD6;
14'd15321:data <=32'hFFFAFFDB;14'd15322:data <=32'hFFF6FFE1;14'd15323:data <=32'hFFF4FFE7;
14'd15324:data <=32'hFFF3FFEF;14'd15325:data <=32'hFFF5FFF5;14'd15326:data <=32'hFFF9FFFC;
14'd15327:data <=32'h00000000;14'd15328:data <=32'h00090002;14'd15329:data <=32'h00120000;
14'd15330:data <=32'h001AFFF9;14'd15331:data <=32'h001FFFEF;14'd15332:data <=32'h001FFFE4;
14'd15333:data <=32'h001BFFD9;14'd15334:data <=32'h0014FFD0;14'd15335:data <=32'h000AFFCB;
14'd15336:data <=32'hFFFFFFC8;14'd15337:data <=32'hFFF5FFC9;14'd15338:data <=32'hFFECFFCD;
14'd15339:data <=32'hFFE5FFD2;14'd15340:data <=32'hFFE0FFD8;14'd15341:data <=32'hFFDDFFDE;
14'd15342:data <=32'hFFDCFFE3;14'd15343:data <=32'hFFDBFFE8;14'd15344:data <=32'hFFDCFFED;
14'd15345:data <=32'hFFDEFFF0;14'd15346:data <=32'hFFE0FFF1;14'd15347:data <=32'hFFE2FFF1;
14'd15348:data <=32'hFFE2FFEE;14'd15349:data <=32'hFFE1FFEB;14'd15350:data <=32'hFFDCFFE7;
14'd15351:data <=32'hFFD3FFE5;14'd15352:data <=32'hFFC8FFE6;14'd15353:data <=32'hFFBDFFEC;
14'd15354:data <=32'hFFB3FFF7;14'd15355:data <=32'hFFAC0005;14'd15356:data <=32'hFFAA0016;
14'd15357:data <=32'hFFAD0026;14'd15358:data <=32'hFFB30035;14'd15359:data <=32'hFFBC0041;
14'd15360:data <=32'hFF9C0023;14'd15361:data <=32'hFF98003F;14'd15362:data <=32'hFFA00052;
14'd15363:data <=32'hFFC8003B;14'd15364:data <=32'hFFEA003F;14'd15365:data <=32'hFFF0003F;
14'd15366:data <=32'hFFF6003F;14'd15367:data <=32'hFFFB003F;14'd15368:data <=32'h0000003E;
14'd15369:data <=32'h0004003D;14'd15370:data <=32'h0007003D;14'd15371:data <=32'h000B0040;
14'd15372:data <=32'h00100043;14'd15373:data <=32'h00190046;14'd15374:data <=32'h00250048;
14'd15375:data <=32'h00340046;14'd15376:data <=32'h0042003E;14'd15377:data <=32'h004F0032;
14'd15378:data <=32'h00580021;14'd15379:data <=32'h005C000F;14'd15380:data <=32'h005BFFFD;
14'd15381:data <=32'h0055FFEC;14'd15382:data <=32'h004BFFDE;14'd15383:data <=32'h003FFFD3;
14'd15384:data <=32'h0032FFCC;14'd15385:data <=32'h0023FFC8;14'd15386:data <=32'h0015FFC8;
14'd15387:data <=32'h0007FFCB;14'd15388:data <=32'hFFFBFFD2;14'd15389:data <=32'hFFF2FFDC;
14'd15390:data <=32'hFFECFFE8;14'd15391:data <=32'hFFECFFF6;14'd15392:data <=32'hFFF00002;
14'd15393:data <=32'hFFF9000C;14'd15394:data <=32'h00040011;14'd15395:data <=32'h00100012;
14'd15396:data <=32'h001B000E;14'd15397:data <=32'h00230006;14'd15398:data <=32'h0028FFFE;
14'd15399:data <=32'h002AFFF5;14'd15400:data <=32'h002AFFED;14'd15401:data <=32'h0028FFE5;
14'd15402:data <=32'h0026FFDF;14'd15403:data <=32'h0023FFD8;14'd15404:data <=32'h001FFFD2;
14'd15405:data <=32'h001BFFCC;14'd15406:data <=32'h0015FFC6;14'd15407:data <=32'h000DFFC1;
14'd15408:data <=32'h0005FFBD;14'd15409:data <=32'hFFFCFFBA;14'd15410:data <=32'hFFF2FFBA;
14'd15411:data <=32'hFFE9FFBB;14'd15412:data <=32'hFFE0FFBC;14'd15413:data <=32'hFFD6FFBE;
14'd15414:data <=32'hFFCCFFC2;14'd15415:data <=32'hFFC1FFC7;14'd15416:data <=32'hFFB7FFCF;
14'd15417:data <=32'hFFADFFDA;14'd15418:data <=32'hFFA6FFE9;14'd15419:data <=32'hFFA2FFFA;
14'd15420:data <=32'hFFA4000C;14'd15421:data <=32'hFFAA001B;14'd15422:data <=32'hFFB50028;
14'd15423:data <=32'hFFC10030;14'd15424:data <=32'hFFACFFD3;14'd15425:data <=32'hFF96FFE3;
14'd15426:data <=32'hFF8EFFFE;14'd15427:data <=32'hFFCA002A;14'd15428:data <=32'hFFEC0029;
14'd15429:data <=32'hFFF00023;14'd15430:data <=32'hFFF1001E;14'd15431:data <=32'hFFF00019;
14'd15432:data <=32'hFFED0016;14'd15433:data <=32'hFFE70015;14'd15434:data <=32'hFFE10017;
14'd15435:data <=32'hFFDB001C;14'd15436:data <=32'hFFD70027;14'd15437:data <=32'hFFD70034;
14'd15438:data <=32'hFFDD0041;14'd15439:data <=32'hFFE9004D;14'd15440:data <=32'hFFF80056;
14'd15441:data <=32'h000A0058;14'd15442:data <=32'h001D0055;14'd15443:data <=32'h002D004D;
14'd15444:data <=32'h00390041;14'd15445:data <=32'h00420034;14'd15446:data <=32'h00470025;
14'd15447:data <=32'h00490017;14'd15448:data <=32'h0048000A;14'd15449:data <=32'h0044FFFD;
14'd15450:data <=32'h003EFFF2;14'd15451:data <=32'h0035FFE8;14'd15452:data <=32'h002AFFE2;
14'd15453:data <=32'h001FFFDF;14'd15454:data <=32'h0013FFDF;14'd15455:data <=32'h0009FFE4;
14'd15456:data <=32'h0002FFEA;14'd15457:data <=32'hFFFEFFF2;14'd15458:data <=32'hFFFEFFF9;
14'd15459:data <=32'hFFFF0000;14'd15460:data <=32'h00020005;14'd15461:data <=32'h00050008;
14'd15462:data <=32'h0008000A;14'd15463:data <=32'h000B000D;14'd15464:data <=32'h000F0010;
14'd15465:data <=32'h00150013;14'd15466:data <=32'h001D0015;14'd15467:data <=32'h00260015;
14'd15468:data <=32'h00310012;14'd15469:data <=32'h003C000A;14'd15470:data <=32'h0046FFFE;
14'd15471:data <=32'h004CFFF0;14'd15472:data <=32'h004EFFDF;14'd15473:data <=32'h004CFFCD;
14'd15474:data <=32'h0046FFBC;14'd15475:data <=32'h003CFFAC;14'd15476:data <=32'h002FFF9F;
14'd15477:data <=32'h001EFF93;14'd15478:data <=32'h000AFF8B;14'd15479:data <=32'hFFF3FF87;
14'd15480:data <=32'hFFDBFF88;14'd15481:data <=32'hFFC3FF90;14'd15482:data <=32'hFFADFF9F;
14'd15483:data <=32'hFF9CFFB3;14'd15484:data <=32'hFF91FFCB;14'd15485:data <=32'hFF8EFFE4;
14'd15486:data <=32'hFF92FFFC;14'd15487:data <=32'hFF9C0010;14'd15488:data <=32'hFFD2FFD1;
14'd15489:data <=32'hFFC3FFD2;14'd15490:data <=32'hFFAEFFDC;14'd15491:data <=32'hFF9F000D;
14'd15492:data <=32'hFFC20017;14'd15493:data <=32'hFFCA001A;14'd15494:data <=32'hFFD1001B;
14'd15495:data <=32'hFFD6001B;14'd15496:data <=32'hFFDA001A;14'd15497:data <=32'hFFDC0018;
14'd15498:data <=32'hFFDB0017;14'd15499:data <=32'hFFDA0017;14'd15500:data <=32'hFFD7001B;
14'd15501:data <=32'hFFD60021;14'd15502:data <=32'hFFD70029;14'd15503:data <=32'hFFDB0031;
14'd15504:data <=32'hFFE30039;14'd15505:data <=32'hFFED003D;14'd15506:data <=32'hFFF8003E;
14'd15507:data <=32'h0002003B;14'd15508:data <=32'h00090037;14'd15509:data <=32'h000F0031;
14'd15510:data <=32'h0012002C;14'd15511:data <=32'h00140028;14'd15512:data <=32'h00160025;
14'd15513:data <=32'h00180022;14'd15514:data <=32'h001B001F;14'd15515:data <=32'h001D001B;
14'd15516:data <=32'h001E0017;14'd15517:data <=32'h001E0013;14'd15518:data <=32'h001D000F;
14'd15519:data <=32'h001C000C;14'd15520:data <=32'h001B000A;14'd15521:data <=32'h001B0008;
14'd15522:data <=32'h001A0005;14'd15523:data <=32'h00190002;14'd15524:data <=32'h0017FFFF;
14'd15525:data <=32'h0014FFFC;14'd15526:data <=32'h000EFFFA;14'd15527:data <=32'h0008FFFB;
14'd15528:data <=32'h0001FFFF;14'd15529:data <=32'hFFFD0007;14'd15530:data <=32'hFFFC0011;
14'd15531:data <=32'hFFFF001C;14'd15532:data <=32'h00070026;14'd15533:data <=32'h0014002D;
14'd15534:data <=32'h0023002F;14'd15535:data <=32'h0033002D;14'd15536:data <=32'h00420025;
14'd15537:data <=32'h00500019;14'd15538:data <=32'h005A000B;14'd15539:data <=32'h0061FFF9;
14'd15540:data <=32'h0064FFE6;14'd15541:data <=32'h0063FFD1;14'd15542:data <=32'h005CFFBC;
14'd15543:data <=32'h0051FFA8;14'd15544:data <=32'h003FFF97;14'd15545:data <=32'h002AFF8B;
14'd15546:data <=32'h0012FF84;14'd15547:data <=32'hFFF9FF85;14'd15548:data <=32'hFFE2FF8C;
14'd15549:data <=32'hFFD0FF98;14'd15550:data <=32'hFFC3FFA7;14'd15551:data <=32'hFFBBFFB7;
14'd15552:data <=32'hFFCBFFC0;14'd15553:data <=32'hFFC1FFC4;14'd15554:data <=32'hFFB7FFC2;
14'd15555:data <=32'hFFB4FFAE;14'd15556:data <=32'hFFC4FFBA;14'd15557:data <=32'hFFBBFFC2;
14'd15558:data <=32'hFFB2FFCC;14'd15559:data <=32'hFFABFFD8;14'd15560:data <=32'hFFA6FFE4;
14'd15561:data <=32'hFFA4FFF2;14'd15562:data <=32'hFFA4FFFF;14'd15563:data <=32'hFFA6000C;
14'd15564:data <=32'hFFA90019;14'd15565:data <=32'hFFAF0027;14'd15566:data <=32'hFFB80033;
14'd15567:data <=32'hFFC4003E;14'd15568:data <=32'hFFD40045;14'd15569:data <=32'hFFE50048;
14'd15570:data <=32'hFFF50044;14'd15571:data <=32'h0003003D;14'd15572:data <=32'h000D0032;
14'd15573:data <=32'h00110025;14'd15574:data <=32'h0011001A;14'd15575:data <=32'h000D0011;
14'd15576:data <=32'h0008000C;14'd15577:data <=32'h0001000A;14'd15578:data <=32'hFFFC000A;
14'd15579:data <=32'hFFF8000C;14'd15580:data <=32'hFFF5000F;14'd15581:data <=32'hFFF40013;
14'd15582:data <=32'hFFF30017;14'd15583:data <=32'hFFF4001C;14'd15584:data <=32'hFFF70021;
14'd15585:data <=32'hFFFC0025;14'd15586:data <=32'h00020027;14'd15587:data <=32'h000A0027;
14'd15588:data <=32'h00100024;14'd15589:data <=32'h0015001F;14'd15590:data <=32'h00170018;
14'd15591:data <=32'h00150012;14'd15592:data <=32'h0012000D;14'd15593:data <=32'h000D000C;
14'd15594:data <=32'h0008000F;14'd15595:data <=32'h00050014;14'd15596:data <=32'h0005001A;
14'd15597:data <=32'h00080021;14'd15598:data <=32'h000F0026;14'd15599:data <=32'h00170029;
14'd15600:data <=32'h00200029;14'd15601:data <=32'h00290027;14'd15602:data <=32'h00310024;
14'd15603:data <=32'h0039001E;14'd15604:data <=32'h00400017;14'd15605:data <=32'h0047000F;
14'd15606:data <=32'h004B0005;14'd15607:data <=32'h004FFFF9;14'd15608:data <=32'h004FFFED;
14'd15609:data <=32'h004DFFE0;14'd15610:data <=32'h0047FFD5;14'd15611:data <=32'h0040FFCB;
14'd15612:data <=32'h0038FFC5;14'd15613:data <=32'h0030FFC0;14'd15614:data <=32'h002AFFBD;
14'd15615:data <=32'h0025FFB9;14'd15616:data <=32'h0003FF96;14'd15617:data <=32'hFFF4FF94;
14'd15618:data <=32'hFFEEFF98;14'd15619:data <=32'h0020FFA2;14'd15620:data <=32'h002DFF9A;
14'd15621:data <=32'h001BFF8E;14'd15622:data <=32'h0006FF86;14'd15623:data <=32'hFFEEFF84;
14'd15624:data <=32'hFFD7FF88;14'd15625:data <=32'hFFC1FF92;14'd15626:data <=32'hFFAEFF9F;
14'd15627:data <=32'hFF9DFFB0;14'd15628:data <=32'hFF91FFC5;14'd15629:data <=32'hFF89FFDC;
14'd15630:data <=32'hFF87FFF5;14'd15631:data <=32'hFF8C000F;14'd15632:data <=32'hFF970026;
14'd15633:data <=32'hFFA90038;14'd15634:data <=32'hFFBE0043;14'd15635:data <=32'hFFD40047;
14'd15636:data <=32'hFFE80044;14'd15637:data <=32'hFFF9003D;14'd15638:data <=32'h00040031;
14'd15639:data <=32'h000B0026;14'd15640:data <=32'h000D001B;14'd15641:data <=32'h000C0011;
14'd15642:data <=32'h00090009;14'd15643:data <=32'h00050003;14'd15644:data <=32'h0000FFFF;
14'd15645:data <=32'hFFFBFFFC;14'd15646:data <=32'hFFF4FFFB;14'd15647:data <=32'hFFEDFFFD;
14'd15648:data <=32'hFFE70000;14'd15649:data <=32'hFFE30005;14'd15650:data <=32'hFFE0000C;
14'd15651:data <=32'hFFE10013;14'd15652:data <=32'hFFE30019;14'd15653:data <=32'hFFE5001D;
14'd15654:data <=32'hFFE90021;14'd15655:data <=32'hFFEB0023;14'd15656:data <=32'hFFEE0026;
14'd15657:data <=32'hFFEF0029;14'd15658:data <=32'hFFF2002E;14'd15659:data <=32'hFFF60033;
14'd15660:data <=32'hFFFC0038;14'd15661:data <=32'h0005003C;14'd15662:data <=32'h000F003E;
14'd15663:data <=32'h001B003C;14'd15664:data <=32'h00250036;14'd15665:data <=32'h002D002F;
14'd15666:data <=32'h00310026;14'd15667:data <=32'h0034001D;14'd15668:data <=32'h00340015;
14'd15669:data <=32'h0032000F;14'd15670:data <=32'h0030000A;14'd15671:data <=32'h002E0006;
14'd15672:data <=32'h002C0004;14'd15673:data <=32'h00290002;14'd15674:data <=32'h00280001;
14'd15675:data <=32'h00260003;14'd15676:data <=32'h00270005;14'd15677:data <=32'h002B0008;
14'd15678:data <=32'h00320009;14'd15679:data <=32'h003C0008;14'd15680:data <=32'h004DFFD1;
14'd15681:data <=32'h004CFFC4;14'd15682:data <=32'h0043FFC1;14'd15683:data <=32'h0044FFED;
14'd15684:data <=32'h0061FFE2;14'd15685:data <=32'h005FFFCC;14'd15686:data <=32'h0056FFB7;
14'd15687:data <=32'h0048FFA6;14'd15688:data <=32'h0037FF98;14'd15689:data <=32'h0023FF8F;
14'd15690:data <=32'h000EFF8A;14'd15691:data <=32'hFFF8FF8A;14'd15692:data <=32'hFFE3FF8E;
14'd15693:data <=32'hFFCFFF97;14'd15694:data <=32'hFFBDFFA5;14'd15695:data <=32'hFFAFFFB7;
14'd15696:data <=32'hFFA7FFCB;14'd15697:data <=32'hFFA5FFE0;14'd15698:data <=32'hFFA9FFF3;
14'd15699:data <=32'hFFB10002;14'd15700:data <=32'hFFBB000E;14'd15701:data <=32'hFFC60014;
14'd15702:data <=32'hFFCF0018;14'd15703:data <=32'hFFD80019;14'd15704:data <=32'hFFDF001A;
14'd15705:data <=32'hFFE5001B;14'd15706:data <=32'hFFEB001B;14'd15707:data <=32'hFFF2001A;
14'd15708:data <=32'hFFF80017;14'd15709:data <=32'hFFFE0012;14'd15710:data <=32'h0001000C;
14'd15711:data <=32'h00030005;14'd15712:data <=32'h0002FFFE;14'd15713:data <=32'hFFFEFFF8;
14'd15714:data <=32'hFFF9FFF4;14'd15715:data <=32'hFFF3FFF1;14'd15716:data <=32'hFFEDFFEF;
14'd15717:data <=32'hFFE5FFEF;14'd15718:data <=32'hFFDEFFF0;14'd15719:data <=32'hFFD5FFF4;
14'd15720:data <=32'hFFCCFFFA;14'd15721:data <=32'hFFC50003;14'd15722:data <=32'hFFBF0010;
14'd15723:data <=32'hFFBD001F;14'd15724:data <=32'hFFBF002F;14'd15725:data <=32'hFFC7003F;
14'd15726:data <=32'hFFD4004D;14'd15727:data <=32'hFFE50056;14'd15728:data <=32'hFFF7005A;
14'd15729:data <=32'h00090058;14'd15730:data <=32'h00180052;14'd15731:data <=32'h00250048;
14'd15732:data <=32'h002D003E;14'd15733:data <=32'h00320033;14'd15734:data <=32'h00340028;
14'd15735:data <=32'h0034001E;14'd15736:data <=32'h00320016;14'd15737:data <=32'h002E0010;
14'd15738:data <=32'h0029000C;14'd15739:data <=32'h0024000A;14'd15740:data <=32'h001F000C;
14'd15741:data <=32'h001D0010;14'd15742:data <=32'h001F0016;14'd15743:data <=32'h0024001C;
14'd15744:data <=32'h00290020;14'd15745:data <=32'h00380022;14'd15746:data <=32'h0040001A;
14'd15747:data <=32'h00340004;14'd15748:data <=32'h00520002;14'd15749:data <=32'h0053FFF4;
14'd15750:data <=32'h0050FFE6;14'd15751:data <=32'h0049FFD9;14'd15752:data <=32'h0042FFCF;
14'd15753:data <=32'h0039FFC8;14'd15754:data <=32'h0030FFC3;14'd15755:data <=32'h0027FFBF;
14'd15756:data <=32'h001DFFBC;14'd15757:data <=32'h0013FFBA;14'd15758:data <=32'h0009FFBB;
14'd15759:data <=32'h0000FFBD;14'd15760:data <=32'hFFF8FFC1;14'd15761:data <=32'hFFF2FFC7;
14'd15762:data <=32'hFFEFFFCC;14'd15763:data <=32'hFFECFFD0;14'd15764:data <=32'hFFEBFFD2;
14'd15765:data <=32'hFFE8FFD3;14'd15766:data <=32'hFFE4FFD4;14'd15767:data <=32'hFFDEFFD6;
14'd15768:data <=32'hFFD6FFDA;14'd15769:data <=32'hFFD1FFE2;14'd15770:data <=32'hFFCCFFEC;
14'd15771:data <=32'hFFCCFFF7;14'd15772:data <=32'hFFCF0001;14'd15773:data <=32'hFFD5000A;
14'd15774:data <=32'hFFDE0010;14'd15775:data <=32'hFFE70013;14'd15776:data <=32'hFFF00012;
14'd15777:data <=32'hFFF90010;14'd15778:data <=32'hFFFF000B;14'd15779:data <=32'h00040003;
14'd15780:data <=32'h0006FFFB;14'd15781:data <=32'h0006FFF2;14'd15782:data <=32'h0003FFE9;
14'd15783:data <=32'hFFFCFFE1;14'd15784:data <=32'hFFF1FFDA;14'd15785:data <=32'hFFE3FFD6;
14'd15786:data <=32'hFFD5FFD8;14'd15787:data <=32'hFFC6FFDF;14'd15788:data <=32'hFFBAFFEA;
14'd15789:data <=32'hFFB2FFFA;14'd15790:data <=32'hFFAF000B;14'd15791:data <=32'hFFB1001C;
14'd15792:data <=32'hFFB7002A;14'd15793:data <=32'hFFC00036;14'd15794:data <=32'hFFCA003E;
14'd15795:data <=32'hFFD50045;14'd15796:data <=32'hFFDF0048;14'd15797:data <=32'hFFE9004B;
14'd15798:data <=32'hFFF2004C;14'd15799:data <=32'hFFFB004D;14'd15800:data <=32'h0004004D;
14'd15801:data <=32'h000D004B;14'd15802:data <=32'h00150048;14'd15803:data <=32'h001C0045;
14'd15804:data <=32'h00220041;14'd15805:data <=32'h0028003E;14'd15806:data <=32'h002E003C;
14'd15807:data <=32'h00360039;14'd15808:data <=32'hFFF90016;14'd15809:data <=32'hFFFD0028;
14'd15810:data <=32'h000E0033;14'd15811:data <=32'h004D0024;14'd15812:data <=32'h006B001A;
14'd15813:data <=32'h006A0004;14'd15814:data <=32'h0064FFF0;14'd15815:data <=32'h0058FFE0;
14'd15816:data <=32'h004AFFD5;14'd15817:data <=32'h003AFFCE;14'd15818:data <=32'h002DFFCD;
14'd15819:data <=32'h0021FFCF;14'd15820:data <=32'h0017FFD3;14'd15821:data <=32'h0011FFD7;
14'd15822:data <=32'h000CFFDD;14'd15823:data <=32'h0009FFE3;14'd15824:data <=32'h0009FFE9;
14'd15825:data <=32'h000BFFEE;14'd15826:data <=32'h0010FFF1;14'd15827:data <=32'h0016FFF0;
14'd15828:data <=32'h001CFFEC;14'd15829:data <=32'h0020FFE4;14'd15830:data <=32'h001FFFDA;
14'd15831:data <=32'h001AFFD1;14'd15832:data <=32'h0012FFC8;14'd15833:data <=32'h0006FFC4;
14'd15834:data <=32'hFFFAFFC4;14'd15835:data <=32'hFFEEFFC8;14'd15836:data <=32'hFFE5FFCF;
14'd15837:data <=32'hFFDFFFD8;14'd15838:data <=32'hFFDCFFE1;14'd15839:data <=32'hFFDCFFEA;
14'd15840:data <=32'hFFDEFFF2;14'd15841:data <=32'hFFE2FFF7;14'd15842:data <=32'hFFE6FFFC;
14'd15843:data <=32'hFFEBFFFF;14'd15844:data <=32'hFFF10001;14'd15845:data <=32'hFFF7FFFF;
14'd15846:data <=32'hFFFCFFFC;14'd15847:data <=32'h0000FFF7;14'd15848:data <=32'h0002FFF0;
14'd15849:data <=32'h0000FFE8;14'd15850:data <=32'hFFFBFFE2;14'd15851:data <=32'hFFF4FFDD;
14'd15852:data <=32'hFFECFFDC;14'd15853:data <=32'hFFE4FFDC;14'd15854:data <=32'hFFDDFFDE;
14'd15855:data <=32'hFFD6FFE2;14'd15856:data <=32'hFFD2FFE6;14'd15857:data <=32'hFFCDFFE9;
14'd15858:data <=32'hFFC8FFEC;14'd15859:data <=32'hFFC3FFF0;14'd15860:data <=32'hFFBBFFF6;
14'd15861:data <=32'hFFB3FFFE;14'd15862:data <=32'hFFAD0009;14'd15863:data <=32'hFFA80018;
14'd15864:data <=32'hFFA70028;14'd15865:data <=32'hFFAB003A;14'd15866:data <=32'hFFB2004B;
14'd15867:data <=32'hFFBD005A;14'd15868:data <=32'hFFCA0067;14'd15869:data <=32'hFFDC0073;
14'd15870:data <=32'hFFEF007B;14'd15871:data <=32'h00040080;14'd15872:data <=32'hFFFC001B;
14'd15873:data <=32'hFFF80029;14'd15874:data <=32'hFFFA003E;14'd15875:data <=32'h00240076;
14'd15876:data <=32'h00540070;14'd15877:data <=32'h00650058;14'd15878:data <=32'h006F003E;
14'd15879:data <=32'h00710023;14'd15880:data <=32'h006B000C;14'd15881:data <=32'h0061FFF9;
14'd15882:data <=32'h0055FFEB;14'd15883:data <=32'h0047FFE2;14'd15884:data <=32'h003AFFDD;
14'd15885:data <=32'h002EFFDB;14'd15886:data <=32'h0023FFDB;14'd15887:data <=32'h0019FFDE;
14'd15888:data <=32'h0012FFE4;14'd15889:data <=32'h000DFFEA;14'd15890:data <=32'h000CFFF2;
14'd15891:data <=32'h000EFFF8;14'd15892:data <=32'h0013FFFB;14'd15893:data <=32'h0019FFFB;
14'd15894:data <=32'h001EFFF7;14'd15895:data <=32'h0021FFF1;14'd15896:data <=32'h0021FFEA;
14'd15897:data <=32'h001EFFE5;14'd15898:data <=32'h0019FFE0;14'd15899:data <=32'h0013FFDF;
14'd15900:data <=32'h000FFFDF;14'd15901:data <=32'h000BFFE0;14'd15902:data <=32'h0009FFE1;
14'd15903:data <=32'h0008FFE1;14'd15904:data <=32'h0007FFE1;14'd15905:data <=32'h0005FFE0;
14'd15906:data <=32'h0002FFDF;14'd15907:data <=32'hFFFFFFDE;14'd15908:data <=32'hFFFCFFDF;
14'd15909:data <=32'hFFF9FFE0;14'd15910:data <=32'hFFF7FFE2;14'd15911:data <=32'hFFF5FFE4;
14'd15912:data <=32'hFFF4FFE6;14'd15913:data <=32'hFFF4FFE7;14'd15914:data <=32'hFFF3FFE8;
14'd15915:data <=32'hFFF2FFEA;14'd15916:data <=32'hFFF1FFEB;14'd15917:data <=32'hFFF2FFEE;
14'd15918:data <=32'hFFF4FFEF;14'd15919:data <=32'hFFF7FFEF;14'd15920:data <=32'hFFFBFFEC;
14'd15921:data <=32'hFFFEFFE7;14'd15922:data <=32'hFFFEFFDE;14'd15923:data <=32'hFFFAFFD4;
14'd15924:data <=32'hFFF1FFCA;14'd15925:data <=32'hFFE4FFC2;14'd15926:data <=32'hFFD2FFC0;
14'd15927:data <=32'hFFBFFFC3;14'd15928:data <=32'hFFADFFCC;14'd15929:data <=32'hFF9DFFDA;
14'd15930:data <=32'hFF90FFEC;14'd15931:data <=32'hFF880001;14'd15932:data <=32'hFF850019;
14'd15933:data <=32'hFF870032;14'd15934:data <=32'hFF8E004A;14'd15935:data <=32'hFF9C0061;
14'd15936:data <=32'hFFC60031;14'd15937:data <=32'hFFC40044;14'd15938:data <=32'hFFC10052;
14'd15939:data <=32'hFFB50069;14'd15940:data <=32'hFFE5007A;14'd15941:data <=32'hFFFC0077;
14'd15942:data <=32'h00100070;14'd15943:data <=32'h00200064;14'd15944:data <=32'h002C0058;
14'd15945:data <=32'h0032004C;14'd15946:data <=32'h00380042;14'd15947:data <=32'h003C0038;
14'd15948:data <=32'h003F002F;14'd15949:data <=32'h00420025;14'd15950:data <=32'h0043001B;
14'd15951:data <=32'h00420011;14'd15952:data <=32'h003F0008;14'd15953:data <=32'h003C0000;
14'd15954:data <=32'h0037FFFB;14'd15955:data <=32'h0033FFF6;14'd15956:data <=32'h002FFFF2;
14'd15957:data <=32'h002CFFEE;14'd15958:data <=32'h0028FFEA;14'd15959:data <=32'h0023FFE6;
14'd15960:data <=32'h001BFFE3;14'd15961:data <=32'h0014FFE3;14'd15962:data <=32'h000BFFE5;
14'd15963:data <=32'h0005FFEA;14'd15964:data <=32'h0001FFF1;14'd15965:data <=32'h0001FFF9;
14'd15966:data <=32'h00050001;14'd15967:data <=32'h000B0005;14'd15968:data <=32'h00130006;
14'd15969:data <=32'h001B0004;14'd15970:data <=32'h0021FFFF;14'd15971:data <=32'h0025FFF8;
14'd15972:data <=32'h0026FFF0;14'd15973:data <=32'h0025FFE9;14'd15974:data <=32'h0022FFE2;
14'd15975:data <=32'h001EFFDC;14'd15976:data <=32'h0018FFD7;14'd15977:data <=32'h0012FFD3;
14'd15978:data <=32'h000BFFD1;14'd15979:data <=32'h0003FFD2;14'd15980:data <=32'hFFFCFFD4;
14'd15981:data <=32'hFFF7FFD8;14'd15982:data <=32'hFFF4FFDF;14'd15983:data <=32'hFFF4FFE4;
14'd15984:data <=32'hFFF7FFE8;14'd15985:data <=32'hFFFDFFEA;14'd15986:data <=32'h0003FFE7;
14'd15987:data <=32'h0006FFE1;14'd15988:data <=32'h0007FFD7;14'd15989:data <=32'h0003FFCD;
14'd15990:data <=32'hFFFAFFC4;14'd15991:data <=32'hFFEEFFBE;14'd15992:data <=32'hFFE0FFBB;
14'd15993:data <=32'hFFD1FFBD;14'd15994:data <=32'hFFC3FFC2;14'd15995:data <=32'hFFB6FFCA;
14'd15996:data <=32'hFFABFFD6;14'd15997:data <=32'hFFA1FFE3;14'd15998:data <=32'hFF9AFFF3;
14'd15999:data <=32'hFF970004;14'd16000:data <=32'hFF8FFFE7;14'd16001:data <=32'hFF7D0000;
14'd16002:data <=32'hFF7B0015;14'd16003:data <=32'hFFA1000F;14'd16004:data <=32'hFFBF0024;
14'd16005:data <=32'hFFC50028;14'd16006:data <=32'hFFCB002C;14'd16007:data <=32'hFFCE002E;
14'd16008:data <=32'hFFD00031;14'd16009:data <=32'hFFD10037;14'd16010:data <=32'hFFD3003F;
14'd16011:data <=32'hFFD90048;14'd16012:data <=32'hFFE20051;14'd16013:data <=32'hFFEF0059;
14'd16014:data <=32'hFFFE005D;14'd16015:data <=32'h000E005C;14'd16016:data <=32'h001E0059;
14'd16017:data <=32'h002C0051;14'd16018:data <=32'h00390047;14'd16019:data <=32'h0043003B;
14'd16020:data <=32'h004A002D;14'd16021:data <=32'h004F001E;14'd16022:data <=32'h0050000D;
14'd16023:data <=32'h004DFFFC;14'd16024:data <=32'h0044FFEC;14'd16025:data <=32'h0038FFE0;
14'd16026:data <=32'h0028FFD9;14'd16027:data <=32'h0018FFD7;14'd16028:data <=32'h0009FFDC;
14'd16029:data <=32'hFFFDFFE4;14'd16030:data <=32'hFFF6FFF0;14'd16031:data <=32'hFFF4FFFC;
14'd16032:data <=32'hFFF70007;14'd16033:data <=32'hFFFD0010;14'd16034:data <=32'h00050015;
14'd16035:data <=32'h000D0018;14'd16036:data <=32'h00140018;14'd16037:data <=32'h001C0016;
14'd16038:data <=32'h00230013;14'd16039:data <=32'h002A000E;14'd16040:data <=32'h00300008;
14'd16041:data <=32'h00340000;14'd16042:data <=32'h0035FFF8;14'd16043:data <=32'h0035FFEF;
14'd16044:data <=32'h0033FFE6;14'd16045:data <=32'h002FFFE0;14'd16046:data <=32'h002AFFDA;
14'd16047:data <=32'h0026FFD6;14'd16048:data <=32'h0023FFD3;14'd16049:data <=32'h0020FFD0;
14'd16050:data <=32'h001DFFCB;14'd16051:data <=32'h001AFFC5;14'd16052:data <=32'h0015FFBE;
14'd16053:data <=32'h000CFFB7;14'd16054:data <=32'h0001FFB2;14'd16055:data <=32'hFFF3FFB0;
14'd16056:data <=32'hFFE5FFB2;14'd16057:data <=32'hFFD8FFB7;14'd16058:data <=32'hFFCEFFC0;
14'd16059:data <=32'hFFC6FFCA;14'd16060:data <=32'hFFC1FFD4;14'd16061:data <=32'hFFBFFFDE;
14'd16062:data <=32'hFFBEFFE7;14'd16063:data <=32'hFFBEFFF0;14'd16064:data <=32'hFFC8FF9D;
14'd16065:data <=32'hFFA9FFA3;14'd16066:data <=32'hFF95FFB9;14'd16067:data <=32'hFFC0FFF6;
14'd16068:data <=32'hFFDD0004;14'd16069:data <=32'hFFE20000;14'd16070:data <=32'hFFE2FFFA;
14'd16071:data <=32'hFFDFFFF4;14'd16072:data <=32'hFFD7FFF0;14'd16073:data <=32'hFFCCFFF0;
14'd16074:data <=32'hFFC0FFF5;14'd16075:data <=32'hFFB60000;14'd16076:data <=32'hFFAF0010;
14'd16077:data <=32'hFFAF0021;14'd16078:data <=32'hFFB30032;14'd16079:data <=32'hFFBC0042;
14'd16080:data <=32'hFFC9004E;14'd16081:data <=32'hFFD90058;14'd16082:data <=32'hFFE9005D;
14'd16083:data <=32'hFFFA005F;14'd16084:data <=32'h000C005D;14'd16085:data <=32'h001D0057;
14'd16086:data <=32'h002D004D;14'd16087:data <=32'h0038003F;14'd16088:data <=32'h0040002E;
14'd16089:data <=32'h0042001C;14'd16090:data <=32'h003F000C;14'd16091:data <=32'h0037FFFE;
14'd16092:data <=32'h002CFFF5;14'd16093:data <=32'h0021FFF0;14'd16094:data <=32'h0016FFEF;
14'd16095:data <=32'h000DFFF2;14'd16096:data <=32'h0007FFF5;14'd16097:data <=32'h0002FFFA;
14'd16098:data <=32'hFFFFFFFE;14'd16099:data <=32'hFFFD0002;14'd16100:data <=32'hFFFB0007;
14'd16101:data <=32'hFFFA000D;14'd16102:data <=32'hFFFA0014;14'd16103:data <=32'hFFFE001C;
14'd16104:data <=32'h00030023;14'd16105:data <=32'h000B0028;14'd16106:data <=32'h0014002C;
14'd16107:data <=32'h0020002D;14'd16108:data <=32'h002B002B;14'd16109:data <=32'h00360027;
14'd16110:data <=32'h00400020;14'd16111:data <=32'h004A0018;14'd16112:data <=32'h0053000D;
14'd16113:data <=32'h005A0000;14'd16114:data <=32'h005FFFEF;14'd16115:data <=32'h0061FFDC;
14'd16116:data <=32'h005EFFC8;14'd16117:data <=32'h0054FFB3;14'd16118:data <=32'h0045FFA1;
14'd16119:data <=32'h0031FF93;14'd16120:data <=32'h0019FF8C;14'd16121:data <=32'h0001FF8C;
14'd16122:data <=32'hFFEBFF91;14'd16123:data <=32'hFFD8FF9D;14'd16124:data <=32'hFFCAFFAB;
14'd16125:data <=32'hFFC1FFBA;14'd16126:data <=32'hFFBCFFCA;14'd16127:data <=32'hFFBBFFD9;
14'd16128:data <=32'h0001FFB3;14'd16129:data <=32'hFFEFFFAA;14'd16130:data <=32'hFFD6FFAB;
14'd16131:data <=32'hFFB5FFDB;14'd16132:data <=32'hFFD2FFF1;14'd16133:data <=32'hFFD8FFF3;
14'd16134:data <=32'hFFDEFFF2;14'd16135:data <=32'hFFE1FFEF;14'd16136:data <=32'hFFE0FFE9;
14'd16137:data <=32'hFFDBFFE6;14'd16138:data <=32'hFFD3FFE5;14'd16139:data <=32'hFFCAFFE9;
14'd16140:data <=32'hFFC2FFF0;14'd16141:data <=32'hFFBDFFFA;14'd16142:data <=32'hFFBB0006;
14'd16143:data <=32'hFFBD0011;14'd16144:data <=32'hFFC0001A;14'd16145:data <=32'hFFC60022;
14'd16146:data <=32'hFFCC002A;14'd16147:data <=32'hFFD30030;14'd16148:data <=32'hFFDA0035;
14'd16149:data <=32'hFFE30038;14'd16150:data <=32'hFFED003A;14'd16151:data <=32'hFFF7003A;
14'd16152:data <=32'h00000036;14'd16153:data <=32'h00070032;14'd16154:data <=32'h000C002B;
14'd16155:data <=32'h000E0025;14'd16156:data <=32'h000F0020;14'd16157:data <=32'h000F001D;
14'd16158:data <=32'h0010001B;14'd16159:data <=32'h00110019;14'd16160:data <=32'h00120017;
14'd16161:data <=32'h00150013;14'd16162:data <=32'h0016000D;14'd16163:data <=32'h00140008;
14'd16164:data <=32'h00100002;14'd16165:data <=32'h0009FFFE;14'd16166:data <=32'h0001FFFD;
14'd16167:data <=32'hFFF9FFFF;14'd16168:data <=32'hFFF20006;14'd16169:data <=32'hFFED000F;
14'd16170:data <=32'hFFEB001A;14'd16171:data <=32'hFFED0025;14'd16172:data <=32'hFFF20030;
14'd16173:data <=32'hFFFB003A;14'd16174:data <=32'h00060042;14'd16175:data <=32'h00140048;
14'd16176:data <=32'h0025004B;14'd16177:data <=32'h00380049;14'd16178:data <=32'h004C0042;
14'd16179:data <=32'h005E0036;14'd16180:data <=32'h006D0023;14'd16181:data <=32'h0077000C;
14'd16182:data <=32'h007BFFF2;14'd16183:data <=32'h0076FFD9;14'd16184:data <=32'h006BFFC2;
14'd16185:data <=32'h005BFFB0;14'd16186:data <=32'h0048FFA3;14'd16187:data <=32'h0035FF9D;
14'd16188:data <=32'h0022FF9A;14'd16189:data <=32'h0011FF9C;14'd16190:data <=32'h0002FF9F;
14'd16191:data <=32'hFFF5FFA4;14'd16192:data <=32'h0001FFB8;14'd16193:data <=32'hFFF8FFB4;
14'd16194:data <=32'hFFEFFFAD;14'd16195:data <=32'hFFEAFF99;14'd16196:data <=32'hFFF5FFAC;
14'd16197:data <=32'hFFEDFFAF;14'd16198:data <=32'hFFE4FFB2;14'd16199:data <=32'hFFDCFFB5;
14'd16200:data <=32'hFFD3FFB9;14'd16201:data <=32'hFFC9FFBE;14'd16202:data <=32'hFFBDFFC6;
14'd16203:data <=32'hFFB5FFD2;14'd16204:data <=32'hFFAEFFE0;14'd16205:data <=32'hFFACFFF0;
14'd16206:data <=32'hFFAF0001;14'd16207:data <=32'hFFB6000F;14'd16208:data <=32'hFFC10019;
14'd16209:data <=32'hFFCC001F;14'd16210:data <=32'hFFD70021;14'd16211:data <=32'hFFE10020;
14'd16212:data <=32'hFFE8001E;14'd16213:data <=32'hFFED001A;14'd16214:data <=32'hFFF10017;
14'd16215:data <=32'hFFF40013;14'd16216:data <=32'hFFF4000F;14'd16217:data <=32'hFFF4000A;
14'd16218:data <=32'hFFF10008;14'd16219:data <=32'hFFED0007;14'd16220:data <=32'hFFE70008;
14'd16221:data <=32'hFFE4000C;14'd16222:data <=32'hFFE10013;14'd16223:data <=32'hFFE3001A;
14'd16224:data <=32'hFFE70021;14'd16225:data <=32'hFFEE0025;14'd16226:data <=32'hFFF60027;
14'd16227:data <=32'hFFFE0024;14'd16228:data <=32'h00040020;14'd16229:data <=32'h00070019;
14'd16230:data <=32'h00060013;14'd16231:data <=32'h0003000E;14'd16232:data <=32'hFFFF000B;
14'd16233:data <=32'hFFF9000B;14'd16234:data <=32'hFFF4000E;14'd16235:data <=32'hFFF00012;
14'd16236:data <=32'hFFEE0018;14'd16237:data <=32'hFFED001F;14'd16238:data <=32'hFFED0027;
14'd16239:data <=32'hFFF0002F;14'd16240:data <=32'hFFF60038;14'd16241:data <=32'hFFFF0040;
14'd16242:data <=32'h000A0046;14'd16243:data <=32'h00190049;14'd16244:data <=32'h00280048;
14'd16245:data <=32'h00370042;14'd16246:data <=32'h00430038;14'd16247:data <=32'h004D002C;
14'd16248:data <=32'h0052001F;14'd16249:data <=32'h00540013;14'd16250:data <=32'h00540008;
14'd16251:data <=32'h0054FFFF;14'd16252:data <=32'h0053FFF6;14'd16253:data <=32'h0054FFEE;
14'd16254:data <=32'h0054FFE4;14'd16255:data <=32'h0053FFD9;14'd16256:data <=32'h0035FFB0;
14'd16257:data <=32'h002AFFA8;14'd16258:data <=32'h0024FFA8;14'd16259:data <=32'h0051FFBD;
14'd16260:data <=32'h005FFFBD;14'd16261:data <=32'h0055FFAB;14'd16262:data <=32'h0047FF9B;
14'd16263:data <=32'h0036FF8E;14'd16264:data <=32'h0021FF84;14'd16265:data <=32'h0008FF7E;
14'd16266:data <=32'hFFEEFF7E;14'd16267:data <=32'hFFD4FF86;14'd16268:data <=32'hFFBDFF95;
14'd16269:data <=32'hFFABFFA9;14'd16270:data <=32'hFFA0FFC1;14'd16271:data <=32'hFF9DFFDA;
14'd16272:data <=32'hFFA1FFF1;14'd16273:data <=32'hFFAA0004;14'd16274:data <=32'hFFB70012;
14'd16275:data <=32'hFFC5001B;14'd16276:data <=32'hFFD20020;14'd16277:data <=32'hFFE00021;
14'd16278:data <=32'hFFEB001F;14'd16279:data <=32'hFFF5001A;14'd16280:data <=32'hFFFD0014;
14'd16281:data <=32'h0002000C;14'd16282:data <=32'h00030002;14'd16283:data <=32'h0001FFF9;
14'd16284:data <=32'hFFFBFFF2;14'd16285:data <=32'hFFF3FFEF;14'd16286:data <=32'hFFEBFFEF;
14'd16287:data <=32'hFFE4FFF2;14'd16288:data <=32'hFFDFFFF7;14'd16289:data <=32'hFFDDFFFD;
14'd16290:data <=32'hFFDC0003;14'd16291:data <=32'hFFDE0007;14'd16292:data <=32'hFFDF0009;
14'd16293:data <=32'hFFE0000B;14'd16294:data <=32'hFFE0000D;14'd16295:data <=32'hFFDE000F;
14'd16296:data <=32'hFFDD0013;14'd16297:data <=32'hFFDC0017;14'd16298:data <=32'hFFDD001D;
14'd16299:data <=32'hFFE00023;14'd16300:data <=32'hFFE30028;14'd16301:data <=32'hFFE9002C;
14'd16302:data <=32'hFFEE002F;14'd16303:data <=32'hFFF30030;14'd16304:data <=32'hFFF80031;
14'd16305:data <=32'hFFFD0032;14'd16306:data <=32'h00030033;14'd16307:data <=32'h00080032;
14'd16308:data <=32'h000D0030;14'd16309:data <=32'h0012002D;14'd16310:data <=32'h00150029;
14'd16311:data <=32'h00170025;14'd16312:data <=32'h00160023;14'd16313:data <=32'h00140023;
14'd16314:data <=32'h00130026;14'd16315:data <=32'h0014002C;14'd16316:data <=32'h00190033;
14'd16317:data <=32'h00220039;14'd16318:data <=32'h0030003C;14'd16319:data <=32'h0040003A;
14'd16320:data <=32'h005C0001;14'd16321:data <=32'h0060FFF5;14'd16322:data <=32'h0059FFEF;
14'd16323:data <=32'h004F001E;14'd16324:data <=32'h006F0020;14'd16325:data <=32'h0078000B;
14'd16326:data <=32'h007CFFF4;14'd16327:data <=32'h007BFFDC;14'd16328:data <=32'h0074FFC4;
14'd16329:data <=32'h0067FFAD;14'd16330:data <=32'h0054FF9A;14'd16331:data <=32'h003CFF8C;
14'd16332:data <=32'h0021FF86;14'd16333:data <=32'h0007FF88;14'd16334:data <=32'hFFF0FF90;
14'd16335:data <=32'hFFDDFF9D;14'd16336:data <=32'hFFD0FFAD;14'd16337:data <=32'hFFC9FFBD;
14'd16338:data <=32'hFFC5FFCC;14'd16339:data <=32'hFFC4FFD9;14'd16340:data <=32'hFFC6FFE5;
14'd16341:data <=32'hFFC9FFF0;14'd16342:data <=32'hFFCDFFF9;14'd16343:data <=32'hFFD30001;
14'd16344:data <=32'hFFDA0007;14'd16345:data <=32'hFFE3000B;14'd16346:data <=32'hFFEB000B;
14'd16347:data <=32'hFFF20009;14'd16348:data <=32'hFFF70006;14'd16349:data <=32'hFFFA0002;
14'd16350:data <=32'hFFFCFFFE;14'd16351:data <=32'hFFFDFFFA;14'd16352:data <=32'hFFFCFFF7;
14'd16353:data <=32'hFFFDFFF4;14'd16354:data <=32'hFFFCFFEF;14'd16355:data <=32'hFFFBFFEB;
14'd16356:data <=32'hFFF8FFE5;14'd16357:data <=32'hFFF1FFDF;14'd16358:data <=32'hFFE8FFDC;
14'd16359:data <=32'hFFDDFFDB;14'd16360:data <=32'hFFD1FFDE;14'd16361:data <=32'hFFC5FFE6;
14'd16362:data <=32'hFFBCFFF1;14'd16363:data <=32'hFFB7FFFF;14'd16364:data <=32'hFFB5000D;
14'd16365:data <=32'hFFB8001C;14'd16366:data <=32'hFFBF0029;14'd16367:data <=32'hFFC70033;
14'd16368:data <=32'hFFD2003B;14'd16369:data <=32'hFFDD0040;14'd16370:data <=32'hFFE80042;
14'd16371:data <=32'hFFF40042;14'd16372:data <=32'hFFFF0040;14'd16373:data <=32'h00080039;
14'd16374:data <=32'h000E0032;14'd16375:data <=32'h00110029;14'd16376:data <=32'h000F0020;
14'd16377:data <=32'h000A001B;14'd16378:data <=32'h00030019;14'd16379:data <=32'hFFFC001D;
14'd16380:data <=32'hFFF80025;14'd16381:data <=32'hFFF80030;14'd16382:data <=32'hFFFD003B;
14'd16383:data <=32'h00070045;
        
        endcase
        
end    
    
    assign dout = data;
    
endmodule
